module drawEnemy(
	input clk,
	input wire [9:0] characterPositionX,
	input wire [8:0] characterPositionY,
	input wire [9:0] drawingPositionX,
	input wire [8:0] drawingPositionY,
	output reg [2:0] rgb
);
	reg [9:0] x;
	reg [9:0] y;
	initial begin
		x = 'd0;
		y = 'd0;
	end

	always @(posedge clk) begin
		x <= (drawingPositionX - characterPositionX + 16);
		y <= (drawingPositionY - characterPositionY + 16);
		if(x==4 && y==1) begin	rgb <= 3'b001;	end
		else if(x==5 && y==1) begin	rgb <= 3'b001;	end
		else if(x==6 && y==1) begin	rgb <= 3'b001;	end
		else if(x==7 && y==1) begin	rgb <= 3'b001;	end
		else if(x==20 && y==1) begin	rgb <= 3'b001;	end
		else if(x==21 && y==1) begin	rgb <= 3'b001;	end
		else if(x==22 && y==1) begin	rgb <= 3'b001;	end
		else if(x==4 && y==2) begin	rgb <= 3'b001;	end
		else if(x==5 && y==2) begin	rgb <= 3'b001;	end
		else if(x==6 && y==2) begin	rgb <= 3'b001;	end
		else if(x==7 && y==2) begin	rgb <= 3'b001;	end
		else if(x==8 && y==2) begin	rgb <= 3'b001;	end
		else if(x==18 && y==2) begin	rgb <= 3'b001;	end
		else if(x==19 && y==2) begin	rgb <= 3'b001;	end
		else if(x==20 && y==2) begin	rgb <= 3'b001;	end
		else if(x==21 && y==2) begin	rgb <= 3'b001;	end
		else if(x==22 && y==2) begin	rgb <= 3'b001;	end
		else if(x==4 && y==3) begin	rgb <= 3'b001;	end
		else if(x==5 && y==3) begin	rgb <= 3'b001;	end
		else if(x==6 && y==3) begin	rgb <= 3'b001;	end
		else if(x==7 && y==3) begin	rgb <= 3'b001;	end
		else if(x==8 && y==3) begin	rgb <= 3'b001;	end
		else if(x==9 && y==3) begin	rgb <= 3'b101;	end
		else if(x==10 && y==3) begin	rgb <= 3'b101;	end
		else if(x==11 && y==3) begin	rgb <= 3'b101;	end
		else if(x==12 && y==3) begin	rgb <= 3'b101;	end
		else if(x==13 && y==3) begin	rgb <= 3'b101;	end
		else if(x==14 && y==3) begin	rgb <= 3'b101;	end
		else if(x==15 && y==3) begin	rgb <= 3'b101;	end
		else if(x==16 && y==3) begin	rgb <= 3'b101;	end
		else if(x==17 && y==3) begin	rgb <= 3'b001;	end
		else if(x==18 && y==3) begin	rgb <= 3'b001;	end
		else if(x==19 && y==3) begin	rgb <= 3'b001;	end
		else if(x==20 && y==3) begin	rgb <= 3'b001;	end
		else if(x==21 && y==3) begin	rgb <= 3'b001;	end
		else if(x==22 && y==3) begin	rgb <= 3'b001;	end
		else if(x==4 && y==4) begin	rgb <= 3'b001;	end
		else if(x==5 && y==4) begin	rgb <= 3'b001;	end
		else if(x==6 && y==4) begin	rgb <= 3'b101;	end
		else if(x==7 && y==4) begin	rgb <= 3'b101;	end
		else if(x==8 && y==4) begin	rgb <= 3'b101;	end
		else if(x==9 && y==4) begin	rgb <= 3'b101;	end
		else if(x==10 && y==4) begin	rgb <= 3'b101;	end
		else if(x==11 && y==4) begin	rgb <= 3'b101;	end
		else if(x==12 && y==4) begin	rgb <= 3'b101;	end
		else if(x==13 && y==4) begin	rgb <= 3'b101;	end
		else if(x==14 && y==4) begin	rgb <= 3'b101;	end
		else if(x==15 && y==4) begin	rgb <= 3'b101;	end
		else if(x==16 && y==4) begin	rgb <= 3'b001;	end
		else if(x==17 && y==4) begin	rgb <= 3'b001;	end
		else if(x==18 && y==4) begin	rgb <= 3'b001;	end
		else if(x==19 && y==4) begin	rgb <= 3'b001;	end
		else if(x==20 && y==4) begin	rgb <= 3'b001;	end
		else if(x==21 && y==4) begin	rgb <= 3'b001;	end
		else if(x==22 && y==4) begin	rgb <= 3'b001;	end
		else if(x==4 && y==5) begin	rgb <= 3'b001;	end
		else if(x==5 && y==5) begin	rgb <= 3'b101;	end
		else if(x==6 && y==5) begin	rgb <= 3'b101;	end
		else if(x==7 && y==5) begin	rgb <= 3'b101;	end
		else if(x==8 && y==5) begin	rgb <= 3'b101;	end
		else if(x==9 && y==5) begin	rgb <= 3'b101;	end
		else if(x==10 && y==5) begin	rgb <= 3'b101;	end
		else if(x==11 && y==5) begin	rgb <= 3'b101;	end
		else if(x==12 && y==5) begin	rgb <= 3'b101;	end
		else if(x==13 && y==5) begin	rgb <= 3'b101;	end
		else if(x==14 && y==5) begin	rgb <= 3'b101;	end
		else if(x==15 && y==5) begin	rgb <= 3'b101;	end
		else if(x==16 && y==5) begin	rgb <= 3'b001;	end
		else if(x==17 && y==5) begin	rgb <= 3'b001;	end
		else if(x==18 && y==5) begin	rgb <= 3'b001;	end
		else if(x==19 && y==5) begin	rgb <= 3'b001;	end
		else if(x==20 && y==5) begin	rgb <= 3'b001;	end
		else if(x==21 && y==5) begin	rgb <= 3'b001;	end
		else if(x==22 && y==5) begin	rgb <= 3'b001;	end
		else if(x==4 && y==6) begin	rgb <= 3'b101;	end
		else if(x==5 && y==6) begin	rgb <= 3'b101;	end
		else if(x==6 && y==6) begin	rgb <= 3'b101;	end
		else if(x==7 && y==6) begin	rgb <= 3'b101;	end
		else if(x==8 && y==6) begin	rgb <= 3'b101;	end
		else if(x==9 && y==6) begin	rgb <= 3'b101;	end
		else if(x==10 && y==6) begin	rgb <= 3'b101;	end
		else if(x==11 && y==6) begin	rgb <= 3'b101;	end
		else if(x==12 && y==6) begin	rgb <= 3'b101;	end
		else if(x==13 && y==6) begin	rgb <= 3'b101;	end
		else if(x==14 && y==6) begin	rgb <= 3'b101;	end
		else if(x==15 && y==6) begin	rgb <= 3'b101;	end
		else if(x==16 && y==6) begin	rgb <= 3'b101;	end
		else if(x==17 && y==6) begin	rgb <= 3'b001;	end
		else if(x==18 && y==6) begin	rgb <= 3'b001;	end
		else if(x==19 && y==6) begin	rgb <= 3'b001;	end
		else if(x==20 && y==6) begin	rgb <= 3'b001;	end
		else if(x==21 && y==6) begin	rgb <= 3'b001;	end
		else if(x==22 && y==6) begin	rgb <= 3'b001;	end
		else if(x==4 && y==7) begin	rgb <= 3'b101;	end
		else if(x==5 && y==7) begin	rgb <= 3'b101;	end
		else if(x==6 && y==7) begin	rgb <= 3'b101;	end
		else if(x==7 && y==7) begin	rgb <= 3'b101;	end
		else if(x==8 && y==7) begin	rgb <= 3'b101;	end
		else if(x==9 && y==7) begin	rgb <= 3'b101;	end
		else if(x==10 && y==7) begin	rgb <= 3'b101;	end
		else if(x==11 && y==7) begin	rgb <= 3'b101;	end
		else if(x==12 && y==7) begin	rgb <= 3'b101;	end
		else if(x==13 && y==7) begin	rgb <= 3'b101;	end
		else if(x==14 && y==7) begin	rgb <= 3'b101;	end
		else if(x==15 && y==7) begin	rgb <= 3'b101;	end
		else if(x==16 && y==7) begin	rgb <= 3'b101;	end
		else if(x==17 && y==7) begin	rgb <= 3'b101;	end
		else if(x==18 && y==7) begin	rgb <= 3'b101;	end
		else if(x==19 && y==7) begin	rgb <= 3'b001;	end
		else if(x==20 && y==7) begin	rgb <= 3'b001;	end
		else if(x==21 && y==7) begin	rgb <= 3'b001;	end
		else if(x==22 && y==7) begin	rgb <= 3'b001;	end
		else if(x==3 && y==8) begin	rgb <= 3'b101;	end
		else if(x==4 && y==8) begin	rgb <= 3'b101;	end
		else if(x==5 && y==8) begin	rgb <= 3'b101;	end
		else if(x==6 && y==8) begin	rgb <= 3'b101;	end
		else if(x==7 && y==8) begin	rgb <= 3'b101;	end
		else if(x==8 && y==8) begin	rgb <= 3'b101;	end
		else if(x==9 && y==8) begin	rgb <= 3'b101;	end
		else if(x==10 && y==8) begin	rgb <= 3'b101;	end
		else if(x==11 && y==8) begin	rgb <= 3'b101;	end
		else if(x==12 && y==8) begin	rgb <= 3'b101;	end
		else if(x==13 && y==8) begin	rgb <= 3'b101;	end
		else if(x==14 && y==8) begin	rgb <= 3'b101;	end
		else if(x==15 && y==8) begin	rgb <= 3'b101;	end
		else if(x==16 && y==8) begin	rgb <= 3'b101;	end
		else if(x==17 && y==8) begin	rgb <= 3'b101;	end
		else if(x==18 && y==8) begin	rgb <= 3'b101;	end
		else if(x==19 && y==8) begin	rgb <= 3'b101;	end
		else if(x==20 && y==8) begin	rgb <= 3'b101;	end
		else if(x==21 && y==8) begin	rgb <= 3'b101;	end
		else if(x==22 && y==8) begin	rgb <= 3'b101;	end
		else if(x==3 && y==9) begin	rgb <= 3'b101;	end
		else if(x==4 && y==9) begin	rgb <= 3'b101;	end
		else if(x==5 && y==9) begin	rgb <= 3'b101;	end
		else if(x==6 && y==9) begin	rgb <= 3'b101;	end
		else if(x==7 && y==9) begin	rgb <= 3'b101;	end
		else if(x==8 && y==9) begin	rgb <= 3'b101;	end
		else if(x==9 && y==9) begin	rgb <= 3'b101;	end
		else if(x==10 && y==9) begin	rgb <= 3'b101;	end
		else if(x==11 && y==9) begin	rgb <= 3'b101;	end
		else if(x==12 && y==9) begin	rgb <= 3'b101;	end
		else if(x==13 && y==9) begin	rgb <= 3'b101;	end
		else if(x==14 && y==9) begin	rgb <= 3'b101;	end
		else if(x==15 && y==9) begin	rgb <= 3'b101;	end
		else if(x==16 && y==9) begin	rgb <= 3'b101;	end
		else if(x==17 && y==9) begin	rgb <= 3'b101;	end
		else if(x==18 && y==9) begin	rgb <= 3'b101;	end
		else if(x==19 && y==9) begin	rgb <= 3'b101;	end
		else if(x==20 && y==9) begin	rgb <= 3'b101;	end
		else if(x==21 && y==9) begin	rgb <= 3'b101;	end
		else if(x==22 && y==9) begin	rgb <= 3'b101;	end
		else if(x==29 && y==9) begin	rgb <= 3'b001;	end
		else if(x==3 && y==10) begin	rgb <= 3'b101;	end
		else if(x==4 && y==10) begin	rgb <= 3'b101;	end
		else if(x==5 && y==10) begin	rgb <= 3'b101;	end
		else if(x==6 && y==10) begin	rgb <= 3'b111;	end
		else if(x==7 && y==10) begin	rgb <= 3'b101;	end
		else if(x==8 && y==10) begin	rgb <= 3'b101;	end
		else if(x==9 && y==10) begin	rgb <= 3'b101;	end
		else if(x==10 && y==10) begin	rgb <= 3'b101;	end
		else if(x==11 && y==10) begin	rgb <= 3'b101;	end
		else if(x==12 && y==10) begin	rgb <= 3'b101;	end
		else if(x==13 && y==10) begin	rgb <= 3'b101;	end
		else if(x==14 && y==10) begin	rgb <= 3'b111;	end
		else if(x==15 && y==10) begin	rgb <= 3'b101;	end
		else if(x==16 && y==10) begin	rgb <= 3'b101;	end
		else if(x==17 && y==10) begin	rgb <= 3'b101;	end
		else if(x==18 && y==10) begin	rgb <= 3'b101;	end
		else if(x==19 && y==10) begin	rgb <= 3'b101;	end
		else if(x==20 && y==10) begin	rgb <= 3'b101;	end
		else if(x==21 && y==10) begin	rgb <= 3'b101;	end
		else if(x==22 && y==10) begin	rgb <= 3'b101;	end
		else if(x==28 && y==10) begin	rgb <= 3'b001;	end
		else if(x==29 && y==10) begin	rgb <= 3'b001;	end
		else if(x==3 && y==11) begin	rgb <= 3'b101;	end
		else if(x==4 && y==11) begin	rgb <= 3'b101;	end
		else if(x==5 && y==11) begin	rgb <= 3'b111;	end
		else if(x==7 && y==11) begin	rgb <= 3'b111;	end
		else if(x==8 && y==11) begin	rgb <= 3'b101;	end
		else if(x==9 && y==11) begin	rgb <= 3'b101;	end
		else if(x==10 && y==11) begin	rgb <= 3'b101;	end
		else if(x==11 && y==11) begin	rgb <= 3'b101;	end
		else if(x==12 && y==11) begin	rgb <= 3'b101;	end
		else if(x==13 && y==11) begin	rgb <= 3'b111;	end
		else if(x==15 && y==11) begin	rgb <= 3'b111;	end
		else if(x==16 && y==11) begin	rgb <= 3'b101;	end
		else if(x==17 && y==11) begin	rgb <= 3'b101;	end
		else if(x==18 && y==11) begin	rgb <= 3'b101;	end
		else if(x==19 && y==11) begin	rgb <= 3'b101;	end
		else if(x==20 && y==11) begin	rgb <= 3'b101;	end
		else if(x==21 && y==11) begin	rgb <= 3'b101;	end
		else if(x==22 && y==11) begin	rgb <= 3'b101;	end
		else if(x==26 && y==11) begin	rgb <= 3'b001;	end
		else if(x==27 && y==11) begin	rgb <= 3'b001;	end
		else if(x==28 && y==11) begin	rgb <= 3'b001;	end
		else if(x==29 && y==11) begin	rgb <= 3'b001;	end
		else if(x==3 && y==12) begin	rgb <= 3'b101;	end
		else if(x==4 && y==12) begin	rgb <= 3'b101;	end
		else if(x==5 && y==12) begin	rgb <= 3'b111;	end
		else if(x==7 && y==12) begin	rgb <= 3'b111;	end
		else if(x==8 && y==12) begin	rgb <= 3'b101;	end
		else if(x==9 && y==12) begin	rgb <= 3'b101;	end
		else if(x==10 && y==12) begin	rgb <= 3'b101;	end
		else if(x==11 && y==12) begin	rgb <= 3'b101;	end
		else if(x==12 && y==12) begin	rgb <= 3'b101;	end
		else if(x==13 && y==12) begin	rgb <= 3'b111;	end
		else if(x==15 && y==12) begin	rgb <= 3'b111;	end
		else if(x==16 && y==12) begin	rgb <= 3'b101;	end
		else if(x==17 && y==12) begin	rgb <= 3'b101;	end
		else if(x==18 && y==12) begin	rgb <= 3'b101;	end
		else if(x==19 && y==12) begin	rgb <= 3'b101;	end
		else if(x==20 && y==12) begin	rgb <= 3'b101;	end
		else if(x==21 && y==12) begin	rgb <= 3'b101;	end
		else if(x==22 && y==12) begin	rgb <= 3'b101;	end
		else if(x==26 && y==12) begin	rgb <= 3'b001;	end
		else if(x==27 && y==12) begin	rgb <= 3'b001;	end
		else if(x==28 && y==12) begin	rgb <= 3'b001;	end
		else if(x==3 && y==13) begin	rgb <= 3'b101;	end
		else if(x==4 && y==13) begin	rgb <= 3'b101;	end
		else if(x==5 && y==13) begin	rgb <= 3'b101;	end
		else if(x==6 && y==13) begin	rgb <= 3'b111;	end
		else if(x==7 && y==13) begin	rgb <= 3'b101;	end
		else if(x==8 && y==13) begin	rgb <= 3'b101;	end
		else if(x==9 && y==13) begin	rgb <= 3'b101;	end
		else if(x==10 && y==13) begin	rgb <= 3'b101;	end
		else if(x==11 && y==13) begin	rgb <= 3'b101;	end
		else if(x==12 && y==13) begin	rgb <= 3'b101;	end
		else if(x==13 && y==13) begin	rgb <= 3'b101;	end
		else if(x==14 && y==13) begin	rgb <= 3'b111;	end
		else if(x==15 && y==13) begin	rgb <= 3'b101;	end
		else if(x==16 && y==13) begin	rgb <= 3'b101;	end
		else if(x==17 && y==13) begin	rgb <= 3'b101;	end
		else if(x==18 && y==13) begin	rgb <= 3'b101;	end
		else if(x==19 && y==13) begin	rgb <= 3'b101;	end
		else if(x==20 && y==13) begin	rgb <= 3'b101;	end
		else if(x==21 && y==13) begin	rgb <= 3'b101;	end
		else if(x==22 && y==13) begin	rgb <= 3'b101;	end
		else if(x==25 && y==13) begin	rgb <= 3'b101;	end
		else if(x==3 && y==14) begin	rgb <= 3'b101;	end
		else if(x==4 && y==14) begin	rgb <= 3'b101;	end
		else if(x==5 && y==14) begin	rgb <= 3'b101;	end
		else if(x==6 && y==14) begin	rgb <= 3'b101;	end
		else if(x==7 && y==14) begin	rgb <= 3'b101;	end
		else if(x==8 && y==14) begin	rgb <= 3'b101;	end
		else if(x==9 && y==14) begin	rgb <= 3'b101;	end
		else if(x==10 && y==14) begin	rgb <= 3'b101;	end
		else if(x==11 && y==14) begin	rgb <= 3'b101;	end
		else if(x==12 && y==14) begin	rgb <= 3'b101;	end
		else if(x==13 && y==14) begin	rgb <= 3'b101;	end
		else if(x==14 && y==14) begin	rgb <= 3'b101;	end
		else if(x==15 && y==14) begin	rgb <= 3'b101;	end
		else if(x==16 && y==14) begin	rgb <= 3'b101;	end
		else if(x==17 && y==14) begin	rgb <= 3'b101;	end
		else if(x==18 && y==14) begin	rgb <= 3'b101;	end
		else if(x==19 && y==14) begin	rgb <= 3'b101;	end
		else if(x==20 && y==14) begin	rgb <= 3'b101;	end
		else if(x==21 && y==14) begin	rgb <= 3'b101;	end
		else if(x==22 && y==14) begin	rgb <= 3'b101;	end
		else if(x==23 && y==14) begin	rgb <= 3'b101;	end
		else if(x==25 && y==14) begin	rgb <= 3'b101;	end
		else if(x==3 && y==15) begin	rgb <= 3'b101;	end
		else if(x==4 && y==15) begin	rgb <= 3'b101;	end
		else if(x==5 && y==15) begin	rgb <= 3'b101;	end
		else if(x==6 && y==15) begin	rgb <= 3'b101;	end
		else if(x==7 && y==15) begin	rgb <= 3'b101;	end
		else if(x==9 && y==15) begin	rgb <= 3'b101;	end
		else if(x==11 && y==15) begin	rgb <= 3'b101;	end
		else if(x==13 && y==15) begin	rgb <= 3'b101;	end
		else if(x==14 && y==15) begin	rgb <= 3'b101;	end
		else if(x==15 && y==15) begin	rgb <= 3'b101;	end
		else if(x==16 && y==15) begin	rgb <= 3'b101;	end
		else if(x==17 && y==15) begin	rgb <= 3'b101;	end
		else if(x==18 && y==15) begin	rgb <= 3'b101;	end
		else if(x==19 && y==15) begin	rgb <= 3'b101;	end
		else if(x==20 && y==15) begin	rgb <= 3'b101;	end
		else if(x==21 && y==15) begin	rgb <= 3'b101;	end
		else if(x==22 && y==15) begin	rgb <= 3'b101;	end
		else if(x==23 && y==15) begin	rgb <= 3'b101;	end
		else if(x==25 && y==15) begin	rgb <= 3'b101;	end
		else if(x==3 && y==16) begin	rgb <= 3'b101;	end
		else if(x==4 && y==16) begin	rgb <= 3'b101;	end
		else if(x==5 && y==16) begin	rgb <= 3'b101;	end
		else if(x==6 && y==16) begin	rgb <= 3'b101;	end
		else if(x==7 && y==16) begin	rgb <= 3'b101;	end
		else if(x==8 && y==16) begin	rgb <= 3'b101;	end
		else if(x==10 && y==16) begin	rgb <= 3'b111;	end
		else if(x==12 && y==16) begin	rgb <= 3'b111;	end
		else if(x==13 && y==16) begin	rgb <= 3'b111;	end
		else if(x==14 && y==16) begin	rgb <= 3'b111;	end
		else if(x==15 && y==16) begin	rgb <= 3'b111;	end
		else if(x==16 && y==16) begin	rgb <= 3'b101;	end
		else if(x==17 && y==16) begin	rgb <= 3'b101;	end
		else if(x==18 && y==16) begin	rgb <= 3'b101;	end
		else if(x==19 && y==16) begin	rgb <= 3'b101;	end
		else if(x==20 && y==16) begin	rgb <= 3'b101;	end
		else if(x==21 && y==16) begin	rgb <= 3'b101;	end
		else if(x==22 && y==16) begin	rgb <= 3'b101;	end
		else if(x==23 && y==16) begin	rgb <= 3'b101;	end
		else if(x==25 && y==16) begin	rgb <= 3'b101;	end
		else if(x==3 && y==17) begin	rgb <= 3'b101;	end
		else if(x==4 && y==17) begin	rgb <= 3'b101;	end
		else if(x==6 && y==17) begin	rgb <= 3'b101;	end
		else if(x==7 && y==17) begin	rgb <= 3'b111;	end
		else if(x==8 && y==17) begin	rgb <= 3'b111;	end
		else if(x==9 && y==17) begin	rgb <= 3'b111;	end
		else if(x==10 && y==17) begin	rgb <= 3'b111;	end
		else if(x==11 && y==17) begin	rgb <= 3'b111;	end
		else if(x==12 && y==17) begin	rgb <= 3'b111;	end
		else if(x==13 && y==17) begin	rgb <= 3'b111;	end
		else if(x==14 && y==17) begin	rgb <= 3'b111;	end
		else if(x==15 && y==17) begin	rgb <= 3'b111;	end
		else if(x==17 && y==17) begin	rgb <= 3'b111;	end
		else if(x==18 && y==17) begin	rgb <= 3'b101;	end
		else if(x==19 && y==17) begin	rgb <= 3'b101;	end
		else if(x==20 && y==17) begin	rgb <= 3'b101;	end
		else if(x==21 && y==17) begin	rgb <= 3'b101;	end
		else if(x==22 && y==17) begin	rgb <= 3'b101;	end
		else if(x==23 && y==17) begin	rgb <= 3'b101;	end
		else if(x==26 && y==17) begin	rgb <= 3'b101;	end
		else if(x==3 && y==18) begin	rgb <= 3'b101;	end
		else if(x==4 && y==18) begin	rgb <= 3'b101;	end
		else if(x==6 && y==18) begin	rgb <= 3'b111;	end
		else if(x==7 && y==18) begin	rgb <= 3'b111;	end
		else if(x==8 && y==18) begin	rgb <= 3'b111;	end
		else if(x==9 && y==18) begin	rgb <= 3'b111;	end
		else if(x==10 && y==18) begin	rgb <= 3'b111;	end
		else if(x==11 && y==18) begin	rgb <= 3'b111;	end
		else if(x==12 && y==18) begin	rgb <= 3'b111;	end
		else if(x==13 && y==18) begin	rgb <= 3'b111;	end
		else if(x==14 && y==18) begin	rgb <= 3'b111;	end
		else if(x==15 && y==18) begin	rgb <= 3'b111;	end
		else if(x==17 && y==18) begin	rgb <= 3'b111;	end
		else if(x==18 && y==18) begin	rgb <= 3'b111;	end
		else if(x==19 && y==18) begin	rgb <= 3'b101;	end
		else if(x==20 && y==18) begin	rgb <= 3'b101;	end
		else if(x==21 && y==18) begin	rgb <= 3'b101;	end
		else if(x==22 && y==18) begin	rgb <= 3'b101;	end
		else if(x==23 && y==18) begin	rgb <= 3'b101;	end
		else if(x==26 && y==18) begin	rgb <= 3'b101;	end
		else if(x==2 && y==19) begin	rgb <= 3'b101;	end
		else if(x==6 && y==19) begin	rgb <= 3'b111;	end
		else if(x==7 && y==19) begin	rgb <= 3'b111;	end
		else if(x==8 && y==19) begin	rgb <= 3'b111;	end
		else if(x==9 && y==19) begin	rgb <= 3'b111;	end
		else if(x==10 && y==19) begin	rgb <= 3'b111;	end
		else if(x==11 && y==19) begin	rgb <= 3'b111;	end
		else if(x==12 && y==19) begin	rgb <= 3'b111;	end
		else if(x==13 && y==19) begin	rgb <= 3'b111;	end
		else if(x==17 && y==19) begin	rgb <= 3'b111;	end
		else if(x==18 && y==19) begin	rgb <= 3'b111;	end
		else if(x==19 && y==19) begin	rgb <= 3'b111;	end
		else if(x==20 && y==19) begin	rgb <= 3'b101;	end
		else if(x==21 && y==19) begin	rgb <= 3'b101;	end
		else if(x==22 && y==19) begin	rgb <= 3'b101;	end
		else if(x==23 && y==19) begin	rgb <= 3'b101;	end
		else if(x==27 && y==19) begin	rgb <= 3'b101;	end
		else if(x==2 && y==20) begin	rgb <= 3'b101;	end
		else if(x==3 && y==20) begin	rgb <= 3'b101;	end
		else if(x==4 && y==20) begin	rgb <= 3'b111;	end
		else if(x==5 && y==20) begin	rgb <= 3'b111;	end
		else if(x==6 && y==20) begin	rgb <= 3'b111;	end
		else if(x==7 && y==20) begin	rgb <= 3'b111;	end
		else if(x==8 && y==20) begin	rgb <= 3'b111;	end
		else if(x==9 && y==20) begin	rgb <= 3'b111;	end
		else if(x==10 && y==20) begin	rgb <= 3'b111;	end
		else if(x==11 && y==20) begin	rgb <= 3'b111;	end
		else if(x==12 && y==20) begin	rgb <= 3'b111;	end
		else if(x==13 && y==20) begin	rgb <= 3'b111;	end
		else if(x==14 && y==20) begin	rgb <= 3'b111;	end
		else if(x==15 && y==20) begin	rgb <= 3'b111;	end
		else if(x==16 && y==20) begin	rgb <= 3'b111;	end
		else if(x==17 && y==20) begin	rgb <= 3'b111;	end
		else if(x==18 && y==20) begin	rgb <= 3'b111;	end
		else if(x==19 && y==20) begin	rgb <= 3'b111;	end
		else if(x==20 && y==20) begin	rgb <= 3'b111;	end
		else if(x==21 && y==20) begin	rgb <= 3'b101;	end
		else if(x==22 && y==20) begin	rgb <= 3'b101;	end
		else if(x==23 && y==20) begin	rgb <= 3'b101;	end
		else if(x==27 && y==20) begin	rgb <= 3'b101;	end
		else if(x==2 && y==21) begin	rgb <= 3'b101;	end
		else if(x==3 && y==21) begin	rgb <= 3'b101;	end
		else if(x==4 && y==21) begin	rgb <= 3'b111;	end
		else if(x==5 && y==21) begin	rgb <= 3'b111;	end
		else if(x==6 && y==21) begin	rgb <= 3'b111;	end
		else if(x==7 && y==21) begin	rgb <= 3'b111;	end
		else if(x==8 && y==21) begin	rgb <= 3'b111;	end
		else if(x==9 && y==21) begin	rgb <= 3'b111;	end
		else if(x==10 && y==21) begin	rgb <= 3'b111;	end
		else if(x==11 && y==21) begin	rgb <= 3'b111;	end
		else if(x==12 && y==21) begin	rgb <= 3'b111;	end
		else if(x==13 && y==21) begin	rgb <= 3'b111;	end
		else if(x==14 && y==21) begin	rgb <= 3'b111;	end
		else if(x==15 && y==21) begin	rgb <= 3'b111;	end
		else if(x==16 && y==21) begin	rgb <= 3'b111;	end
		else if(x==17 && y==21) begin	rgb <= 3'b111;	end
		else if(x==18 && y==21) begin	rgb <= 3'b111;	end
		else if(x==19 && y==21) begin	rgb <= 3'b111;	end
		else if(x==20 && y==21) begin	rgb <= 3'b111;	end
		else if(x==21 && y==21) begin	rgb <= 3'b101;	end
		else if(x==22 && y==21) begin	rgb <= 3'b101;	end
		else if(x==23 && y==21) begin	rgb <= 3'b101;	end
		else if(x==27 && y==21) begin	rgb <= 3'b101;	end
		else if(x==2 && y==22) begin	rgb <= 3'b101;	end
		else if(x==3 && y==22) begin	rgb <= 3'b101;	end
		else if(x==4 && y==22) begin	rgb <= 3'b111;	end
		else if(x==5 && y==22) begin	rgb <= 3'b111;	end
		else if(x==6 && y==22) begin	rgb <= 3'b111;	end
		else if(x==7 && y==22) begin	rgb <= 3'b111;	end
		else if(x==8 && y==22) begin	rgb <= 3'b111;	end
		else if(x==9 && y==22) begin	rgb <= 3'b111;	end
		else if(x==10 && y==22) begin	rgb <= 3'b111;	end
		else if(x==11 && y==22) begin	rgb <= 3'b111;	end
		else if(x==12 && y==22) begin	rgb <= 3'b111;	end
		else if(x==13 && y==22) begin	rgb <= 3'b111;	end
		else if(x==14 && y==22) begin	rgb <= 3'b111;	end
		else if(x==15 && y==22) begin	rgb <= 3'b111;	end
		else if(x==16 && y==22) begin	rgb <= 3'b111;	end
		else if(x==17 && y==22) begin	rgb <= 3'b111;	end
		else if(x==18 && y==22) begin	rgb <= 3'b111;	end
		else if(x==19 && y==22) begin	rgb <= 3'b111;	end
		else if(x==20 && y==22) begin	rgb <= 3'b111;	end
		else if(x==21 && y==22) begin	rgb <= 3'b101;	end
		else if(x==22 && y==22) begin	rgb <= 3'b101;	end
		else if(x==23 && y==22) begin	rgb <= 3'b101;	end
		else if(x==26 && y==22) begin	rgb <= 3'b101;	end
		else if(x==2 && y==23) begin	rgb <= 3'b101;	end
		else if(x==3 && y==23) begin	rgb <= 3'b101;	end
		else if(x==4 && y==23) begin	rgb <= 3'b111;	end
		else if(x==5 && y==23) begin	rgb <= 3'b111;	end
		else if(x==6 && y==23) begin	rgb <= 3'b111;	end
		else if(x==7 && y==23) begin	rgb <= 3'b111;	end
		else if(x==8 && y==23) begin	rgb <= 3'b111;	end
		else if(x==9 && y==23) begin	rgb <= 3'b111;	end
		else if(x==10 && y==23) begin	rgb <= 3'b111;	end
		else if(x==11 && y==23) begin	rgb <= 3'b111;	end
		else if(x==12 && y==23) begin	rgb <= 3'b111;	end
		else if(x==13 && y==23) begin	rgb <= 3'b111;	end
		else if(x==14 && y==23) begin	rgb <= 3'b111;	end
		else if(x==15 && y==23) begin	rgb <= 3'b111;	end
		else if(x==16 && y==23) begin	rgb <= 3'b111;	end
		else if(x==17 && y==23) begin	rgb <= 3'b111;	end
		else if(x==18 && y==23) begin	rgb <= 3'b111;	end
		else if(x==19 && y==23) begin	rgb <= 3'b111;	end
		else if(x==20 && y==23) begin	rgb <= 3'b111;	end
		else if(x==21 && y==23) begin	rgb <= 3'b101;	end
		else if(x==22 && y==23) begin	rgb <= 3'b101;	end
		else if(x==23 && y==23) begin	rgb <= 3'b101;	end
		else if(x==26 && y==23) begin	rgb <= 3'b101;	end
		else if(x==2 && y==24) begin	rgb <= 3'b101;	end
		else if(x==3 && y==24) begin	rgb <= 3'b101;	end
		else if(x==4 && y==24) begin	rgb <= 3'b101;	end
		else if(x==5 && y==24) begin	rgb <= 3'b111;	end
		else if(x==6 && y==24) begin	rgb <= 3'b111;	end
		else if(x==7 && y==24) begin	rgb <= 3'b111;	end
		else if(x==8 && y==24) begin	rgb <= 3'b111;	end
		else if(x==9 && y==24) begin	rgb <= 3'b111;	end
		else if(x==10 && y==24) begin	rgb <= 3'b111;	end
		else if(x==11 && y==24) begin	rgb <= 3'b111;	end
		else if(x==12 && y==24) begin	rgb <= 3'b111;	end
		else if(x==13 && y==24) begin	rgb <= 3'b111;	end
		else if(x==14 && y==24) begin	rgb <= 3'b111;	end
		else if(x==15 && y==24) begin	rgb <= 3'b111;	end
		else if(x==16 && y==24) begin	rgb <= 3'b111;	end
		else if(x==17 && y==24) begin	rgb <= 3'b111;	end
		else if(x==18 && y==24) begin	rgb <= 3'b111;	end
		else if(x==19 && y==24) begin	rgb <= 3'b111;	end
		else if(x==20 && y==24) begin	rgb <= 3'b101;	end
		else if(x==21 && y==24) begin	rgb <= 3'b101;	end
		else if(x==22 && y==24) begin	rgb <= 3'b101;	end
		else if(x==23 && y==24) begin	rgb <= 3'b101;	end
		else if(x==24 && y==24) begin	rgb <= 3'b101;	end
		else if(x==25 && y==24) begin	rgb <= 3'b101;	end
		else if(x==2 && y==25) begin	rgb <= 3'b101;	end
		else if(x==3 && y==25) begin	rgb <= 3'b101;	end
		else if(x==4 && y==25) begin	rgb <= 3'b101;	end
		else if(x==5 && y==25) begin	rgb <= 3'b101;	end
		else if(x==6 && y==25) begin	rgb <= 3'b111;	end
		else if(x==7 && y==25) begin	rgb <= 3'b111;	end
		else if(x==8 && y==25) begin	rgb <= 3'b111;	end
		else if(x==9 && y==25) begin	rgb <= 3'b111;	end
		else if(x==10 && y==25) begin	rgb <= 3'b111;	end
		else if(x==11 && y==25) begin	rgb <= 3'b111;	end
		else if(x==12 && y==25) begin	rgb <= 3'b111;	end
		else if(x==13 && y==25) begin	rgb <= 3'b111;	end
		else if(x==14 && y==25) begin	rgb <= 3'b111;	end
		else if(x==15 && y==25) begin	rgb <= 3'b111;	end
		else if(x==16 && y==25) begin	rgb <= 3'b111;	end
		else if(x==17 && y==25) begin	rgb <= 3'b111;	end
		else if(x==18 && y==25) begin	rgb <= 3'b111;	end
		else if(x==19 && y==25) begin	rgb <= 3'b101;	end
		else if(x==20 && y==25) begin	rgb <= 3'b101;	end
		else if(x==21 && y==25) begin	rgb <= 3'b101;	end
		else if(x==22 && y==25) begin	rgb <= 3'b101;	end
		else if(x==2 && y==26) begin	rgb <= 3'b101;	end
		else if(x==3 && y==26) begin	rgb <= 3'b101;	end
		else if(x==4 && y==26) begin	rgb <= 3'b101;	end
		else if(x==5 && y==26) begin	rgb <= 3'b101;	end
		else if(x==6 && y==26) begin	rgb <= 3'b101;	end
		else if(x==7 && y==26) begin	rgb <= 3'b111;	end
		else if(x==8 && y==26) begin	rgb <= 3'b111;	end
		else if(x==9 && y==26) begin	rgb <= 3'b111;	end
		else if(x==10 && y==26) begin	rgb <= 3'b111;	end
		else if(x==11 && y==26) begin	rgb <= 3'b111;	end
		else if(x==12 && y==26) begin	rgb <= 3'b111;	end
		else if(x==13 && y==26) begin	rgb <= 3'b111;	end
		else if(x==14 && y==26) begin	rgb <= 3'b111;	end
		else if(x==15 && y==26) begin	rgb <= 3'b111;	end
		else if(x==16 && y==26) begin	rgb <= 3'b111;	end
		else if(x==17 && y==26) begin	rgb <= 3'b111;	end
		else if(x==18 && y==26) begin	rgb <= 3'b101;	end
		else if(x==19 && y==26) begin	rgb <= 3'b101;	end
		else if(x==5 && y==27) begin	rgb <= 3'b101;	end
		else if(x==6 && y==27) begin	rgb <= 3'b101;	end
		else if(x==7 && y==27) begin	rgb <= 3'b101;	end
		else if(x==8 && y==27) begin	rgb <= 3'b101;	end
		else if(x==9 && y==27) begin	rgb <= 3'b111;	end
		else if(x==10 && y==27) begin	rgb <= 3'b111;	end
		else if(x==11 && y==27) begin	rgb <= 3'b111;	end
		else if(x==12 && y==27) begin	rgb <= 3'b111;	end
		else if(x==13 && y==27) begin	rgb <= 3'b111;	end
		else if(x==14 && y==27) begin	rgb <= 3'b111;	end
		else if(x==15 && y==27) begin	rgb <= 3'b111;	end
		else if(x==16 && y==27) begin	rgb <= 3'b101;	end
		else if(x==17 && y==27) begin	rgb <= 3'b101;	end
		else if(x==7 && y==28) begin	rgb <= 3'b101;	end
		else if(x==8 && y==28) begin	rgb <= 3'b101;	end
		else if(x==9 && y==28) begin	rgb <= 3'b101;	end
		else if(x==10 && y==28) begin	rgb <= 3'b101;	end
		else if(x==11 && y==28) begin	rgb <= 3'b101;	end
		else if(x==12 && y==28) begin	rgb <= 3'b101;	end
		else if(x==13 && y==28) begin	rgb <= 3'b101;	end
		else if(x==14 && y==28) begin	rgb <= 3'b101;	end
		else if(x==15 && y==28) begin	rgb <= 3'b101;	end
		else begin rgb <= 3'b000; end// Width: 30, Height: 30 From: C:/Users/ITPCC/OneDrive/Documents/CPE223/Gun/pink_beam.png
	end
endmodule
