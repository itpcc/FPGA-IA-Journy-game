module drawMainCharacter(
	input clk,
	input wire [9:0] characterPositionX,
	input wire [8:0] characterPositionY,
	input wire [9:0] drawingPositionX,
	input wire [8:0] drawingPositionY,
	output reg [2:0] rgb
);
	reg [9:0] x;
	reg [9:0] y;
	initial begin
		x = 'd0;
		y = 'd0;
	end

	always @(posedge clk) begin
		x <= (drawingPositionX - characterPositionX + 26);
		y <= (drawingPositionY - characterPositionY + 26);
		if(x == 25 && y == 25 || x == 25 && y == 24 || x == 25 && y == 26 || x == 24 && y == 25 || x == 24 && y == 24 || x == 24 && y == 26 || x == 26 && y == 25 || x == 26 && y == 24 || x == 26 && y == 26 )	begin/*	rgb <= 3'b010;*/	end
		else if(x==27 && y==1) begin	rgb <= 3'b101;	end
		else if(x==28 && y==1) begin	rgb <= 3'b101;	end
		else if(x==29 && y==1) begin	rgb <= 3'b101;	end
		else if(x==30 && y==1) begin	rgb <= 3'b101;	end
		else if(x==31 && y==1) begin	rgb <= 3'b101;	end
		else if(x==25 && y==2) begin	rgb <= 3'b101;	end
		else if(x==26 && y==2) begin	rgb <= 3'b101;	end
		else if(x==27 && y==2) begin	rgb <= 3'b101;	end
		else if(x==28 && y==2) begin	rgb <= 3'b101;	end
		else if(x==29 && y==2) begin	rgb <= 3'b101;	end
		else if(x==25 && y==3) begin	rgb <= 3'b101;	end
		else if(x==26 && y==3) begin	rgb <= 3'b101;	end
		else if(x==27 && y==3) begin	rgb <= 3'b101;	end
		else if(x==28 && y==3) begin	rgb <= 3'b101;	end
		else if(x==29 && y==3) begin	rgb <= 3'b101;	end
		else if(x==25 && y==4) begin	rgb <= 3'b101;	end
		else if(x==26 && y==4) begin	rgb <= 3'b101;	end
		else if(x==27 && y==4) begin	rgb <= 3'b101;	end
		else if(x==28 && y==4) begin	rgb <= 3'b101;	end
		else if(x==29 && y==4) begin	rgb <= 3'b101;	end
		else if(x==22 && y==5) begin	rgb <= 3'b101;	end
		else if(x==23 && y==5) begin	rgb <= 3'b101;	end
		else if(x==24 && y==5) begin	rgb <= 3'b101;	end
		else if(x==25 && y==5) begin	rgb <= 3'b101;	end
		else if(x==26 && y==5) begin	rgb <= 3'b101;	end
		else if(x==22 && y==6) begin	rgb <= 3'b101;	end
		else if(x==23 && y==6) begin	rgb <= 3'b101;	end
		else if(x==24 && y==6) begin	rgb <= 3'b101;	end
		else if(x==25 && y==6) begin	rgb <= 3'b101;	end
		else if(x==26 && y==6) begin	rgb <= 3'b101;	end
		else if(x==17 && y==7) begin	rgb <= 3'b101;	end
		else if(x==18 && y==7) begin	rgb <= 3'b101;	end
		else if(x==19 && y==7) begin	rgb <= 3'b101;	end
		else if(x==20 && y==7) begin	rgb <= 3'b101;	end
		else if(x==21 && y==7) begin	rgb <= 3'b101;	end
		else if(x==22 && y==7) begin	rgb <= 3'b111;	end
		else if(x==23 && y==7) begin	rgb <= 3'b111;	end
		else if(x==24 && y==7) begin	rgb <= 3'b111;	end
		else if(x==25 && y==7) begin	rgb <= 3'b111;	end
		else if(x==26 && y==7) begin	rgb <= 3'b111;	end
		else if(x==27 && y==7) begin	rgb <= 3'b111;	end
		else if(x==28 && y==7) begin	rgb <= 3'b101;	end
		else if(x==29 && y==7) begin	rgb <= 3'b101;	end
		else if(x==30 && y==7) begin	rgb <= 3'b101;	end
		else if(x==31 && y==7) begin	rgb <= 3'b101;	end
		else if(x==17 && y==8) begin	rgb <= 3'b101;	end
		else if(x==18 && y==8) begin	rgb <= 3'b101;	end
		else if(x==19 && y==8) begin	rgb <= 3'b101;	end
		else if(x==20 && y==8) begin	rgb <= 3'b101;	end
		else if(x==21 && y==8) begin	rgb <= 3'b101;	end
		else if(x==22 && y==8) begin	rgb <= 3'b111;	end
		else if(x==23 && y==8) begin	rgb <= 3'b111;	end
		else if(x==24 && y==8) begin	rgb <= 3'b111;	end
		else if(x==25 && y==8) begin	rgb <= 3'b111;	end
		else if(x==26 && y==8) begin	rgb <= 3'b111;	end
		else if(x==27 && y==8) begin	rgb <= 3'b111;	end
		else if(x==28 && y==8) begin	rgb <= 3'b101;	end
		else if(x==29 && y==8) begin	rgb <= 3'b101;	end
		else if(x==30 && y==8) begin	rgb <= 3'b101;	end
		else if(x==31 && y==8) begin	rgb <= 3'b101;	end
		else if(x==12 && y==9) begin	rgb <= 3'b101;	end
		else if(x==13 && y==9) begin	rgb <= 3'b101;	end
		else if(x==14 && y==9) begin	rgb <= 3'b101;	end
		else if(x==15 && y==9) begin	rgb <= 3'b101;	end
		else if(x==16 && y==9) begin	rgb <= 3'b101;	end
		else if(x==17 && y==9) begin	rgb <= 3'b111;	end
		else if(x==18 && y==9) begin	rgb <= 3'b111;	end
		else if(x==19 && y==9) begin	rgb <= 3'b111;	end
		else if(x==20 && y==9) begin	rgb <= 3'b111;	end
		else if(x==21 && y==9) begin	rgb <= 3'b111;	end
		else if(x==22 && y==9) begin	rgb <= 3'b111;	end
		else if(x==23 && y==9) begin	rgb <= 3'b111;	end
		else if(x==24 && y==9) begin	rgb <= 3'b111;	end
		else if(x==25 && y==9) begin	rgb <= 3'b111;	end
		else if(x==26 && y==9) begin	rgb <= 3'b111;	end
		else if(x==27 && y==9) begin	rgb <= 3'b111;	end
		else if(x==28 && y==9) begin	rgb <= 3'b111;	end
		else if(x==29 && y==9) begin	rgb <= 3'b111;	end
		else if(x==30 && y==9) begin	rgb <= 3'b111;	end
		else if(x==31 && y==9) begin	rgb <= 3'b111;	end
		else if(x==32 && y==9) begin	rgb <= 3'b111;	end
		else if(x==33 && y==9) begin	rgb <= 3'b101;	end
		else if(x==34 && y==9) begin	rgb <= 3'b101;	end
		else if(x==35 && y==9) begin	rgb <= 3'b101;	end
		else if(x==36 && y==9) begin	rgb <= 3'b101;	end
		else if(x==37 && y==9) begin	rgb <= 3'b101;	end
		else if(x==12 && y==10) begin	rgb <= 3'b101;	end
		else if(x==13 && y==10) begin	rgb <= 3'b101;	end
		else if(x==14 && y==10) begin	rgb <= 3'b101;	end
		else if(x==15 && y==10) begin	rgb <= 3'b101;	end
		else if(x==16 && y==10) begin	rgb <= 3'b101;	end
		else if(x==17 && y==10) begin	rgb <= 3'b111;	end
		else if(x==18 && y==10) begin	rgb <= 3'b111;	end
		else if(x==19 && y==10) begin	rgb <= 3'b111;	end
		else if(x==20 && y==10) begin	rgb <= 3'b111;	end
		else if(x==21 && y==10) begin	rgb <= 3'b111;	end
		else if(x==22 && y==10) begin	rgb <= 3'b111;	end
		else if(x==23 && y==10) begin	rgb <= 3'b111;	end
		else if(x==24 && y==10) begin	rgb <= 3'b111;	end
		else if(x==25 && y==10) begin	rgb <= 3'b111;	end
		else if(x==26 && y==10) begin	rgb <= 3'b111;	end
		else if(x==27 && y==10) begin	rgb <= 3'b111;	end
		else if(x==28 && y==10) begin	rgb <= 3'b111;	end
		else if(x==29 && y==10) begin	rgb <= 3'b111;	end
		else if(x==30 && y==10) begin	rgb <= 3'b111;	end
		else if(x==31 && y==10) begin	rgb <= 3'b111;	end
		else if(x==32 && y==10) begin	rgb <= 3'b111;	end
		else if(x==33 && y==10) begin	rgb <= 3'b101;	end
		else if(x==34 && y==10) begin	rgb <= 3'b101;	end
		else if(x==35 && y==10) begin	rgb <= 3'b101;	end
		else if(x==36 && y==10) begin	rgb <= 3'b101;	end
		else if(x==10 && y==11) begin	rgb <= 3'b101;	end
		else if(x==11 && y==11) begin	rgb <= 3'b101;	end
		else if(x==12 && y==11) begin	rgb <= 3'b111;	end
		else if(x==13 && y==11) begin	rgb <= 3'b111;	end
		else if(x==14 && y==11) begin	rgb <= 3'b111;	end
		else if(x==15 && y==11) begin	rgb <= 3'b111;	end
		else if(x==16 && y==11) begin	rgb <= 3'b111;	end
		else if(x==17 && y==11) begin	rgb <= 3'b111;	end
		else if(x==18 && y==11) begin	rgb <= 3'b111;	end
		else if(x==19 && y==11) begin	rgb <= 3'b111;	end
		else if(x==20 && y==11) begin	rgb <= 3'b111;	end
		else if(x==21 && y==11) begin	rgb <= 3'b111;	end
		else if(x==22 && y==11) begin	rgb <= 3'b111;	end
		else if(x==23 && y==11) begin	rgb <= 3'b111;	end
		else if(x==24 && y==11) begin	rgb <= 3'b111;	end
		else if(x==25 && y==11) begin	rgb <= 3'b111;	end
		else if(x==26 && y==11) begin	rgb <= 3'b111;	end
		else if(x==27 && y==11) begin	rgb <= 3'b111;	end
		else if(x==28 && y==11) begin	rgb <= 3'b111;	end
		else if(x==29 && y==11) begin	rgb <= 3'b111;	end
		else if(x==30 && y==11) begin	rgb <= 3'b111;	end
		else if(x==31 && y==11) begin	rgb <= 3'b111;	end
		else if(x==32 && y==11) begin	rgb <= 3'b111;	end
		else if(x==33 && y==11) begin	rgb <= 3'b111;	end
		else if(x==34 && y==11) begin	rgb <= 3'b111;	end
		else if(x==35 && y==11) begin	rgb <= 3'b111;	end
		else if(x==36 && y==11) begin	rgb <= 3'b111;	end
		else if(x==37 && y==11) begin	rgb <= 3'b111;	end
		else if(x==38 && y==11) begin	rgb <= 3'b101;	end
		else if(x==39 && y==11) begin	rgb <= 3'b101;	end
		else if(x==10 && y==12) begin	rgb <= 3'b101;	end
		else if(x==11 && y==12) begin	rgb <= 3'b101;	end
		else if(x==12 && y==12) begin	rgb <= 3'b111;	end
		else if(x==13 && y==12) begin	rgb <= 3'b111;	end
		else if(x==14 && y==12) begin	rgb <= 3'b111;	end
		else if(x==15 && y==12) begin	rgb <= 3'b111;	end
		else if(x==16 && y==12) begin	rgb <= 3'b111;	end
		else if(x==17 && y==12) begin	rgb <= 3'b111;	end
		else if(x==18 && y==12) begin	rgb <= 3'b111;	end
		else if(x==19 && y==12) begin	rgb <= 3'b111;	end
		else if(x==20 && y==12) begin	rgb <= 3'b111;	end
		else if(x==21 && y==12) begin	rgb <= 3'b111;	end
		else if(x==22 && y==12) begin	rgb <= 3'b111;	end
		else if(x==23 && y==12) begin	rgb <= 3'b111;	end
		else if(x==24 && y==12) begin	rgb <= 3'b111;	end
		else if(x==25 && y==12) begin	rgb <= 3'b111;	end
		else if(x==26 && y==12) begin	rgb <= 3'b111;	end
		else if(x==27 && y==12) begin	rgb <= 3'b111;	end
		else if(x==28 && y==12) begin	rgb <= 3'b111;	end
		else if(x==29 && y==12) begin	rgb <= 3'b111;	end
		else if(x==30 && y==12) begin	rgb <= 3'b111;	end
		else if(x==31 && y==12) begin	rgb <= 3'b111;	end
		else if(x==32 && y==12) begin	rgb <= 3'b111;	end
		else if(x==33 && y==12) begin	rgb <= 3'b111;	end
		else if(x==34 && y==12) begin	rgb <= 3'b111;	end
		else if(x==35 && y==12) begin	rgb <= 3'b111;	end
		else if(x==36 && y==12) begin	rgb <= 3'b111;	end
		else if(x==37 && y==12) begin	rgb <= 3'b111;	end
		else if(x==38 && y==12) begin	rgb <= 3'b101;	end
		else if(x==39 && y==12) begin	rgb <= 3'b101;	end
		else if(x==10 && y==13) begin	rgb <= 3'b101;	end
		else if(x==11 && y==13) begin	rgb <= 3'b101;	end
		else if(x==12 && y==13) begin	rgb <= 3'b111;	end
		else if(x==13 && y==13) begin	rgb <= 3'b111;	end
		else if(x==14 && y==13) begin	rgb <= 3'b111;	end
		else if(x==15 && y==13) begin	rgb <= 3'b111;	end
		else if(x==16 && y==13) begin	rgb <= 3'b111;	end
		else if(x==17 && y==13) begin	rgb <= 3'b111;	end
		else if(x==18 && y==13) begin	rgb <= 3'b111;	end
		else if(x==19 && y==13) begin	rgb <= 3'b111;	end
		else if(x==20 && y==13) begin	rgb <= 3'b111;	end
		else if(x==21 && y==13) begin	rgb <= 3'b111;	end
		else if(x==22 && y==13) begin	rgb <= 3'b111;	end
		else if(x==23 && y==13) begin	rgb <= 3'b111;	end
		else if(x==24 && y==13) begin	rgb <= 3'b111;	end
		else if(x==25 && y==13) begin	rgb <= 3'b111;	end
		else if(x==26 && y==13) begin	rgb <= 3'b111;	end
		else if(x==27 && y==13) begin	rgb <= 3'b111;	end
		else if(x==28 && y==13) begin	rgb <= 3'b111;	end
		else if(x==29 && y==13) begin	rgb <= 3'b111;	end
		else if(x==30 && y==13) begin	rgb <= 3'b111;	end
		else if(x==31 && y==13) begin	rgb <= 3'b111;	end
		else if(x==32 && y==13) begin	rgb <= 3'b111;	end
		else if(x==33 && y==13) begin	rgb <= 3'b111;	end
		else if(x==34 && y==13) begin	rgb <= 3'b111;	end
		else if(x==35 && y==13) begin	rgb <= 3'b111;	end
		else if(x==36 && y==13) begin	rgb <= 3'b111;	end
		else if(x==37 && y==13) begin	rgb <= 3'b111;	end
		else if(x==38 && y==13) begin	rgb <= 3'b101;	end
		else if(x==39 && y==13) begin	rgb <= 3'b101;	end
		else if(x==7 && y==14) begin	rgb <= 3'b101;	end
		else if(x==8 && y==14) begin	rgb <= 3'b101;	end
		else if(x==9 && y==14) begin	rgb <= 3'b101;	end
		else if(x==10 && y==14) begin	rgb <= 3'b111;	end
		else if(x==11 && y==14) begin	rgb <= 3'b111;	end
		else if(x==12 && y==14) begin	rgb <= 3'b111;	end
		else if(x==13 && y==14) begin	rgb <= 3'b111;	end
		else if(x==14 && y==14) begin	rgb <= 3'b111;	end
		else if(x==15 && y==14) begin	rgb <= 3'b111;	end
		else if(x==16 && y==14) begin	rgb <= 3'b111;	end
		else if(x==17 && y==14) begin	rgb <= 3'b111;	end
		else if(x==18 && y==14) begin	rgb <= 3'b111;	end
		else if(x==19 && y==14) begin	rgb <= 3'b111;	end
		else if(x==20 && y==14) begin	rgb <= 3'b111;	end
		else if(x==21 && y==14) begin	rgb <= 3'b111;	end
		else if(x==22 && y==14) begin	rgb <= 3'b111;	end
		else if(x==23 && y==14) begin	rgb <= 3'b111;	end
		else if(x==24 && y==14) begin	rgb <= 3'b111;	end
		else if(x==25 && y==14) begin	rgb <= 3'b111;	end
		else if(x==26 && y==14) begin	rgb <= 3'b111;	end
		else if(x==27 && y==14) begin	rgb <= 3'b111;	end
		else if(x==28 && y==14) begin	rgb <= 3'b111;	end
		else if(x==29 && y==14) begin	rgb <= 3'b111;	end
		else if(x==30 && y==14) begin	rgb <= 3'b111;	end
		else if(x==31 && y==14) begin	rgb <= 3'b111;	end
		else if(x==32 && y==14) begin	rgb <= 3'b111;	end
		else if(x==33 && y==14) begin	rgb <= 3'b111;	end
		else if(x==34 && y==14) begin	rgb <= 3'b111;	end
		else if(x==35 && y==14) begin	rgb <= 3'b111;	end
		else if(x==36 && y==14) begin	rgb <= 3'b111;	end
		else if(x==37 && y==14) begin	rgb <= 3'b111;	end
		else if(x==38 && y==14) begin	rgb <= 3'b111;	end
		else if(x==39 && y==14) begin	rgb <= 3'b111;	end
		else if(x==40 && y==14) begin	rgb <= 3'b101;	end
		else if(x==41 && y==14) begin	rgb <= 3'b101;	end
		else if(x==7 && y==15) begin	rgb <= 3'b101;	end
		else if(x==8 && y==15) begin	rgb <= 3'b101;	end
		else if(x==9 && y==15) begin	rgb <= 3'b101;	end
		else if(x==10 && y==15) begin	rgb <= 3'b111;	end
		else if(x==11 && y==15) begin	rgb <= 3'b111;	end
		else if(x==12 && y==15) begin	rgb <= 3'b111;	end
		else if(x==13 && y==15) begin	rgb <= 3'b111;	end
		else if(x==14 && y==15) begin	rgb <= 3'b111;	end
		else if(x==15 && y==15) begin	rgb <= 3'b111;	end
		else if(x==16 && y==15) begin	rgb <= 3'b111;	end
		else if(x==17 && y==15) begin	rgb <= 3'b111;	end
		else if(x==18 && y==15) begin	rgb <= 3'b111;	end
		else if(x==19 && y==15) begin	rgb <= 3'b111;	end
		else if(x==20 && y==15) begin	rgb <= 3'b111;	end
		else if(x==21 && y==15) begin	rgb <= 3'b111;	end
		else if(x==22 && y==15) begin	rgb <= 3'b111;	end
		else if(x==23 && y==15) begin	rgb <= 3'b111;	end
		else if(x==24 && y==15) begin	rgb <= 3'b111;	end
		else if(x==25 && y==15) begin	rgb <= 3'b111;	end
		else if(x==26 && y==15) begin	rgb <= 3'b111;	end
		else if(x==27 && y==15) begin	rgb <= 3'b111;	end
		else if(x==28 && y==15) begin	rgb <= 3'b111;	end
		else if(x==29 && y==15) begin	rgb <= 3'b111;	end
		else if(x==30 && y==15) begin	rgb <= 3'b111;	end
		else if(x==31 && y==15) begin	rgb <= 3'b111;	end
		else if(x==32 && y==15) begin	rgb <= 3'b111;	end
		else if(x==33 && y==15) begin	rgb <= 3'b111;	end
		else if(x==34 && y==15) begin	rgb <= 3'b111;	end
		else if(x==35 && y==15) begin	rgb <= 3'b111;	end
		else if(x==36 && y==15) begin	rgb <= 3'b111;	end
		else if(x==37 && y==15) begin	rgb <= 3'b111;	end
		else if(x==38 && y==15) begin	rgb <= 3'b111;	end
		else if(x==39 && y==15) begin	rgb <= 3'b111;	end
		else if(x==40 && y==15) begin	rgb <= 3'b101;	end
		else if(x==41 && y==15) begin	rgb <= 3'b101;	end
		else if(x==7 && y==16) begin	rgb <= 3'b101;	end
		else if(x==8 && y==16) begin	rgb <= 3'b101;	end
		else if(x==9 && y==16) begin	rgb <= 3'b101;	end
		else if(x==10 && y==16) begin	rgb <= 3'b111;	end
		else if(x==11 && y==16) begin	rgb <= 3'b111;	end
		else if(x==12 && y==16) begin	rgb <= 3'b111;	end
		else if(x==13 && y==16) begin	rgb <= 3'b111;	end
		else if(x==14 && y==16) begin	rgb <= 3'b111;	end
		else if(x==15 && y==16) begin	rgb <= 3'b111;	end
		else if(x==16 && y==16) begin	rgb <= 3'b111;	end
		else if(x==17 && y==16) begin	rgb <= 3'b111;	end
		else if(x==18 && y==16) begin	rgb <= 3'b111;	end
		else if(x==19 && y==16) begin	rgb <= 3'b111;	end
		else if(x==20 && y==16) begin	rgb <= 3'b101;	end
		else if(x==21 && y==16) begin	rgb <= 3'b101;	end
		else if(x==22 && y==16) begin	rgb <= 3'b111;	end
		else if(x==23 && y==16) begin	rgb <= 3'b111;	end
		else if(x==24 && y==16) begin	rgb <= 3'b111;	end
		else if(x==25 && y==16) begin	rgb <= 3'b111;	end
		else if(x==26 && y==16) begin	rgb <= 3'b111;	end
		else if(x==27 && y==16) begin	rgb <= 3'b111;	end
		else if(x==28 && y==16) begin	rgb <= 3'b101;	end
		else if(x==29 && y==16) begin	rgb <= 3'b101;	end
		else if(x==30 && y==16) begin	rgb <= 3'b111;	end
		else if(x==31 && y==16) begin	rgb <= 3'b111;	end
		else if(x==32 && y==16) begin	rgb <= 3'b111;	end
		else if(x==33 && y==16) begin	rgb <= 3'b111;	end
		else if(x==34 && y==16) begin	rgb <= 3'b111;	end
		else if(x==35 && y==16) begin	rgb <= 3'b111;	end
		else if(x==36 && y==16) begin	rgb <= 3'b111;	end
		else if(x==37 && y==16) begin	rgb <= 3'b111;	end
		else if(x==38 && y==16) begin	rgb <= 3'b111;	end
		else if(x==39 && y==16) begin	rgb <= 3'b111;	end
		else if(x==40 && y==16) begin	rgb <= 3'b101;	end
		else if(x==41 && y==16) begin	rgb <= 3'b101;	end
		else if(x==7 && y==17) begin	rgb <= 3'b101;	end
		else if(x==8 && y==17) begin	rgb <= 3'b101;	end
		else if(x==9 && y==17) begin	rgb <= 3'b101;	end
		else if(x==10 && y==17) begin	rgb <= 3'b111;	end
		else if(x==11 && y==17) begin	rgb <= 3'b111;	end
		else if(x==12 && y==17) begin	rgb <= 3'b111;	end
		else if(x==13 && y==17) begin	rgb <= 3'b111;	end
		else if(x==14 && y==17) begin	rgb <= 3'b111;	end
		else if(x==15 && y==17) begin	rgb <= 3'b111;	end
		else if(x==16 && y==17) begin	rgb <= 3'b111;	end
		else if(x==17 && y==17) begin	rgb <= 3'b111;	end
		else if(x==18 && y==17) begin	rgb <= 3'b111;	end
		else if(x==19 && y==17) begin	rgb <= 3'b111;	end
		else if(x==20 && y==17) begin	rgb <= 3'b101;	end
		else if(x==21 && y==17) begin	rgb <= 3'b101;	end
		else if(x==22 && y==17) begin	rgb <= 3'b111;	end
		else if(x==23 && y==17) begin	rgb <= 3'b111;	end
		else if(x==24 && y==17) begin	rgb <= 3'b111;	end
		else if(x==25 && y==17) begin	rgb <= 3'b111;	end
		else if(x==26 && y==17) begin	rgb <= 3'b111;	end
		else if(x==27 && y==17) begin	rgb <= 3'b111;	end
		else if(x==28 && y==17) begin	rgb <= 3'b101;	end
		else if(x==29 && y==17) begin	rgb <= 3'b101;	end
		else if(x==30 && y==17) begin	rgb <= 3'b111;	end
		else if(x==31 && y==17) begin	rgb <= 3'b111;	end
		else if(x==32 && y==17) begin	rgb <= 3'b111;	end
		else if(x==33 && y==17) begin	rgb <= 3'b111;	end
		else if(x==34 && y==17) begin	rgb <= 3'b111;	end
		else if(x==35 && y==17) begin	rgb <= 3'b111;	end
		else if(x==36 && y==17) begin	rgb <= 3'b111;	end
		else if(x==37 && y==17) begin	rgb <= 3'b111;	end
		else if(x==38 && y==17) begin	rgb <= 3'b111;	end
		else if(x==39 && y==17) begin	rgb <= 3'b111;	end
		else if(x==40 && y==17) begin	rgb <= 3'b101;	end
		else if(x==41 && y==17) begin	rgb <= 3'b101;	end
		else if(x==5 && y==18) begin	rgb <= 3'b101;	end
		else if(x==6 && y==18) begin	rgb <= 3'b101;	end
		else if(x==7 && y==18) begin	rgb <= 3'b111;	end
		else if(x==8 && y==18) begin	rgb <= 3'b111;	end
		else if(x==9 && y==18) begin	rgb <= 3'b111;	end
		else if(x==10 && y==18) begin	rgb <= 3'b111;	end
		else if(x==11 && y==18) begin	rgb <= 3'b111;	end
		else if(x==12 && y==18) begin	rgb <= 3'b111;	end
		else if(x==13 && y==18) begin	rgb <= 3'b111;	end
		else if(x==14 && y==18) begin	rgb <= 3'b111;	end
		else if(x==15 && y==18) begin	rgb <= 3'b111;	end
		else if(x==16 && y==18) begin	rgb <= 3'b111;	end
		else if(x==17 && y==18) begin	rgb <= 3'b111;	end
		else if(x==18 && y==18) begin	rgb <= 3'b111;	end
		else if(x==19 && y==18) begin	rgb <= 3'b111;	end
		else if(x==20 && y==18) begin	rgb <= 3'b101;	end
		else if(x==21 && y==18) begin	rgb <= 3'b101;	end
		else if(x==22 && y==18) begin	rgb <= 3'b111;	end
		else if(x==23 && y==18) begin	rgb <= 3'b111;	end
		else if(x==24 && y==18) begin	rgb <= 3'b111;	end
		else if(x==25 && y==18) begin	rgb <= 3'b111;	end
		else if(x==26 && y==18) begin	rgb <= 3'b111;	end
		else if(x==27 && y==18) begin	rgb <= 3'b111;	end
		else if(x==28 && y==18) begin	rgb <= 3'b101;	end
		else if(x==29 && y==18) begin	rgb <= 3'b101;	end
		else if(x==30 && y==18) begin	rgb <= 3'b101;	end
		else if(x==31 && y==18) begin	rgb <= 3'b101;	end
		else if(x==32 && y==18) begin	rgb <= 3'b111;	end
		else if(x==33 && y==18) begin	rgb <= 3'b111;	end
		else if(x==34 && y==18) begin	rgb <= 3'b111;	end
		else if(x==35 && y==18) begin	rgb <= 3'b111;	end
		else if(x==36 && y==18) begin	rgb <= 3'b111;	end
		else if(x==37 && y==18) begin	rgb <= 3'b111;	end
		else if(x==38 && y==18) begin	rgb <= 3'b111;	end
		else if(x==39 && y==18) begin	rgb <= 3'b111;	end
		else if(x==40 && y==18) begin	rgb <= 3'b111;	end
		else if(x==41 && y==18) begin	rgb <= 3'b111;	end
		else if(x==42 && y==18) begin	rgb <= 3'b111;	end
		else if(x==43 && y==18) begin	rgb <= 3'b101;	end
		else if(x==44 && y==18) begin	rgb <= 3'b101;	end
		else if(x==5 && y==19) begin	rgb <= 3'b101;	end
		else if(x==6 && y==19) begin	rgb <= 3'b101;	end
		else if(x==7 && y==19) begin	rgb <= 3'b111;	end
		else if(x==8 && y==19) begin	rgb <= 3'b111;	end
		else if(x==9 && y==19) begin	rgb <= 3'b111;	end
		else if(x==10 && y==19) begin	rgb <= 3'b111;	end
		else if(x==11 && y==19) begin	rgb <= 3'b111;	end
		else if(x==12 && y==19) begin	rgb <= 3'b111;	end
		else if(x==13 && y==19) begin	rgb <= 3'b111;	end
		else if(x==14 && y==19) begin	rgb <= 3'b111;	end
		else if(x==15 && y==19) begin	rgb <= 3'b111;	end
		else if(x==16 && y==19) begin	rgb <= 3'b111;	end
		else if(x==17 && y==19) begin	rgb <= 3'b111;	end
		else if(x==18 && y==19) begin	rgb <= 3'b111;	end
		else if(x==19 && y==19) begin	rgb <= 3'b111;	end
		else if(x==20 && y==19) begin	rgb <= 3'b101;	end
		else if(x==21 && y==19) begin	rgb <= 3'b101;	end
		else if(x==22 && y==19) begin	rgb <= 3'b111;	end
		else if(x==23 && y==19) begin	rgb <= 3'b111;	end
		else if(x==24 && y==19) begin	rgb <= 3'b111;	end
		else if(x==25 && y==19) begin	rgb <= 3'b111;	end
		else if(x==26 && y==19) begin	rgb <= 3'b111;	end
		else if(x==27 && y==19) begin	rgb <= 3'b111;	end
		else if(x==28 && y==19) begin	rgb <= 3'b101;	end
		else if(x==29 && y==19) begin	rgb <= 3'b101;	end
		else if(x==30 && y==19) begin	rgb <= 3'b101;	end
		else if(x==31 && y==19) begin	rgb <= 3'b101;	end
		else if(x==32 && y==19) begin	rgb <= 3'b111;	end
		else if(x==33 && y==19) begin	rgb <= 3'b111;	end
		else if(x==34 && y==19) begin	rgb <= 3'b111;	end
		else if(x==35 && y==19) begin	rgb <= 3'b111;	end
		else if(x==36 && y==19) begin	rgb <= 3'b111;	end
		else if(x==37 && y==19) begin	rgb <= 3'b111;	end
		else if(x==38 && y==19) begin	rgb <= 3'b111;	end
		else if(x==39 && y==19) begin	rgb <= 3'b111;	end
		else if(x==40 && y==19) begin	rgb <= 3'b111;	end
		else if(x==41 && y==19) begin	rgb <= 3'b111;	end
		else if(x==42 && y==19) begin	rgb <= 3'b111;	end
		else if(x==43 && y==19) begin	rgb <= 3'b101;	end
		else if(x==44 && y==19) begin	rgb <= 3'b101;	end
		else if(x==5 && y==20) begin	rgb <= 3'b101;	end
		else if(x==6 && y==20) begin	rgb <= 3'b101;	end
		else if(x==7 && y==20) begin	rgb <= 3'b111;	end
		else if(x==8 && y==20) begin	rgb <= 3'b111;	end
		else if(x==9 && y==20) begin	rgb <= 3'b111;	end
		else if(x==10 && y==20) begin	rgb <= 3'b111;	end
		else if(x==11 && y==20) begin	rgb <= 3'b111;	end
		else if(x==12 && y==20) begin	rgb <= 3'b111;	end
		else if(x==13 && y==20) begin	rgb <= 3'b111;	end
		else if(x==14 && y==20) begin	rgb <= 3'b111;	end
		else if(x==15 && y==20) begin	rgb <= 3'b111;	end
		else if(x==16 && y==20) begin	rgb <= 3'b111;	end
		else if(x==17 && y==20) begin	rgb <= 3'b111;	end
		else if(x==18 && y==20) begin	rgb <= 3'b101;	end
		else if(x==19 && y==20) begin	rgb <= 3'b101;	end
		else if(x==20 && y==20) begin	rgb <= 3'b111;	end
		else if(x==21 && y==20) begin	rgb <= 3'b111;	end
		else if(x==22 && y==20) begin	rgb <= 3'b111;	end
		else if(x==23 && y==20) begin	rgb <= 3'b101;	end
		else if(x==24 && y==20) begin	rgb <= 3'b101;	end
		else if(x==25 && y==20) begin	rgb <= 3'b111;	end
		else if(x==26 && y==20) begin	rgb <= 3'b111;	end
		else if(x==27 && y==20) begin	rgb <= 3'b111;	end
		else if(x==28 && y==20) begin	rgb <= 3'b101;	end
		else if(x==29 && y==20) begin	rgb <= 3'b101;	end
		else if(x==30 && y==20) begin	rgb <= 3'b111;	end
		else if(x==31 && y==20) begin	rgb <= 3'b111;	end
		else if(x==32 && y==20) begin	rgb <= 3'b111;	end
		else if(x==33 && y==20) begin	rgb <= 3'b101;	end
		else if(x==34 && y==20) begin	rgb <= 3'b101;	end
		else if(x==35 && y==20) begin	rgb <= 3'b111;	end
		else if(x==36 && y==20) begin	rgb <= 3'b111;	end
		else if(x==37 && y==20) begin	rgb <= 3'b111;	end
		else if(x==38 && y==20) begin	rgb <= 3'b111;	end
		else if(x==39 && y==20) begin	rgb <= 3'b111;	end
		else if(x==40 && y==20) begin	rgb <= 3'b111;	end
		else if(x==41 && y==20) begin	rgb <= 3'b111;	end
		else if(x==42 && y==20) begin	rgb <= 3'b111;	end
		else if(x==43 && y==20) begin	rgb <= 3'b101;	end
		else if(x==44 && y==20) begin	rgb <= 3'b101;	end
		else if(x==5 && y==21) begin	rgb <= 3'b101;	end
		else if(x==6 && y==21) begin	rgb <= 3'b101;	end
		else if(x==7 && y==21) begin	rgb <= 3'b111;	end
		else if(x==8 && y==21) begin	rgb <= 3'b111;	end
		else if(x==9 && y==21) begin	rgb <= 3'b111;	end
		else if(x==10 && y==21) begin	rgb <= 3'b111;	end
		else if(x==11 && y==21) begin	rgb <= 3'b111;	end
		else if(x==12 && y==21) begin	rgb <= 3'b111;	end
		else if(x==13 && y==21) begin	rgb <= 3'b111;	end
		else if(x==14 && y==21) begin	rgb <= 3'b111;	end
		else if(x==15 && y==21) begin	rgb <= 3'b111;	end
		else if(x==16 && y==21) begin	rgb <= 3'b111;	end
		else if(x==17 && y==21) begin	rgb <= 3'b111;	end
		else if(x==18 && y==21) begin	rgb <= 3'b101;	end
		else if(x==19 && y==21) begin	rgb <= 3'b101;	end
		else if(x==20 && y==21) begin	rgb <= 3'b111;	end
		else if(x==21 && y==21) begin	rgb <= 3'b111;	end
		else if(x==22 && y==21) begin	rgb <= 3'b111;	end
		else if(x==23 && y==21) begin	rgb <= 3'b101;	end
		else if(x==24 && y==21) begin	rgb <= 3'b101;	end
		else if(x==25 && y==21) begin	rgb <= 3'b111;	end
		else if(x==26 && y==21) begin	rgb <= 3'b111;	end
		else if(x==27 && y==21) begin	rgb <= 3'b111;	end
		else if(x==28 && y==21) begin	rgb <= 3'b101;	end
		else if(x==29 && y==21) begin	rgb <= 3'b101;	end
		else if(x==30 && y==21) begin	rgb <= 3'b111;	end
		else if(x==31 && y==21) begin	rgb <= 3'b111;	end
		else if(x==32 && y==21) begin	rgb <= 3'b111;	end
		else if(x==33 && y==21) begin	rgb <= 3'b101;	end
		else if(x==34 && y==21) begin	rgb <= 3'b101;	end
		else if(x==35 && y==21) begin	rgb <= 3'b111;	end
		else if(x==36 && y==21) begin	rgb <= 3'b111;	end
		else if(x==37 && y==21) begin	rgb <= 3'b111;	end
		else if(x==38 && y==21) begin	rgb <= 3'b111;	end
		else if(x==39 && y==21) begin	rgb <= 3'b111;	end
		else if(x==40 && y==21) begin	rgb <= 3'b111;	end
		else if(x==41 && y==21) begin	rgb <= 3'b111;	end
		else if(x==42 && y==21) begin	rgb <= 3'b111;	end
		else if(x==43 && y==21) begin	rgb <= 3'b101;	end
		else if(x==44 && y==21) begin	rgb <= 3'b101;	end
		else if(x==5 && y==22) begin	rgb <= 3'b101;	end
		else if(x==6 && y==22) begin	rgb <= 3'b101;	end
		else if(x==7 && y==22) begin	rgb <= 3'b111;	end
		else if(x==8 && y==22) begin	rgb <= 3'b111;	end
		else if(x==9 && y==22) begin	rgb <= 3'b111;	end
		else if(x==10 && y==22) begin	rgb <= 3'b111;	end
		else if(x==11 && y==22) begin	rgb <= 3'b111;	end
		else if(x==12 && y==22) begin	rgb <= 3'b111;	end
		else if(x==13 && y==22) begin	rgb <= 3'b111;	end
		else if(x==14 && y==22) begin	rgb <= 3'b111;	end
		else if(x==15 && y==22) begin	rgb <= 3'b111;	end
		else if(x==16 && y==22) begin	rgb <= 3'b111;	end
		else if(x==17 && y==22) begin	rgb <= 3'b111;	end
		else if(x==18 && y==22) begin	rgb <= 3'b101;	end
		else if(x==19 && y==22) begin	rgb <= 3'b101;	end
		else if(x==20 && y==22) begin	rgb <= 3'b111;	end
		else if(x==21 && y==22) begin	rgb <= 3'b111;	end
		else if(x==22 && y==22) begin	rgb <= 3'b111;	end
		else if(x==23 && y==22) begin	rgb <= 3'b101;	end
		else if(x==24 && y==22) begin	rgb <= 3'b101;	end
		else if(x==25 && y==22) begin	rgb <= 3'b111;	end
		else if(x==26 && y==22) begin	rgb <= 3'b111;	end
		else if(x==27 && y==22) begin	rgb <= 3'b111;	end
		else if(x==28 && y==22) begin	rgb <= 3'b101;	end
		else if(x==29 && y==22) begin	rgb <= 3'b101;	end
		else if(x==30 && y==22) begin	rgb <= 3'b111;	end
		else if(x==31 && y==22) begin	rgb <= 3'b111;	end
		else if(x==32 && y==22) begin	rgb <= 3'b111;	end
		else if(x==33 && y==22) begin	rgb <= 3'b101;	end
		else if(x==34 && y==22) begin	rgb <= 3'b101;	end
		else if(x==35 && y==22) begin	rgb <= 3'b111;	end
		else if(x==36 && y==22) begin	rgb <= 3'b111;	end
		else if(x==37 && y==22) begin	rgb <= 3'b111;	end
		else if(x==38 && y==22) begin	rgb <= 3'b111;	end
		else if(x==39 && y==22) begin	rgb <= 3'b111;	end
		else if(x==40 && y==22) begin	rgb <= 3'b111;	end
		else if(x==41 && y==22) begin	rgb <= 3'b111;	end
		else if(x==42 && y==22) begin	rgb <= 3'b111;	end
		else if(x==43 && y==22) begin	rgb <= 3'b101;	end
		else if(x==44 && y==22) begin	rgb <= 3'b101;	end
		else if(x==5 && y==23) begin	rgb <= 3'b101;	end
		else if(x==6 && y==23) begin	rgb <= 3'b101;	end
		else if(x==7 && y==23) begin	rgb <= 3'b111;	end
		else if(x==8 && y==23) begin	rgb <= 3'b111;	end
		else if(x==9 && y==23) begin	rgb <= 3'b111;	end
		else if(x==10 && y==23) begin	rgb <= 3'b111;	end
		else if(x==11 && y==23) begin	rgb <= 3'b111;	end
		else if(x==12 && y==23) begin	rgb <= 3'b111;	end
		else if(x==13 && y==23) begin	rgb <= 3'b111;	end
		else if(x==14 && y==23) begin	rgb <= 3'b111;	end
		else if(x==15 && y==23) begin	rgb <= 3'b101;	end
		else if(x==16 && y==23) begin	rgb <= 3'b101;	end
		else if(x==17 && y==23) begin	rgb <= 3'b111;	end
		else if(x==18 && y==23) begin	rgb <= 3'b111;	end
		else if(x==19 && y==23) begin	rgb <= 3'b111;	end
		else if(x==20 && y==23) begin	rgb <= 3'b111;	end
		else if(x==21 && y==23) begin	rgb <= 3'b111;	end
		else if(x==22 && y==23) begin	rgb <= 3'b111;	end
		else if(x==23 && y==23) begin	rgb <= 3'b101;	end
		else if(x==24 && y==23) begin	rgb <= 3'b101;	end
		else if(x==25 && y==23) begin	rgb <= 3'b111;	end
		else if(x==26 && y==23) begin	rgb <= 3'b111;	end
		else if(x==27 && y==23) begin	rgb <= 3'b111;	end
		else if(x==28 && y==23) begin	rgb <= 3'b101;	end
		else if(x==29 && y==23) begin	rgb <= 3'b101;	end
		else if(x==30 && y==23) begin	rgb <= 3'b111;	end
		else if(x==31 && y==23) begin	rgb <= 3'b111;	end
		else if(x==32 && y==23) begin	rgb <= 3'b111;	end
		else if(x==33 && y==23) begin	rgb <= 3'b101;	end
		else if(x==34 && y==23) begin	rgb <= 3'b101;	end
		else if(x==35 && y==23) begin	rgb <= 3'b111;	end
		else if(x==36 && y==23) begin	rgb <= 3'b111;	end
		else if(x==37 && y==23) begin	rgb <= 3'b111;	end
		else if(x==38 && y==23) begin	rgb <= 3'b111;	end
		else if(x==39 && y==23) begin	rgb <= 3'b111;	end
		else if(x==40 && y==23) begin	rgb <= 3'b111;	end
		else if(x==41 && y==23) begin	rgb <= 3'b111;	end
		else if(x==42 && y==23) begin	rgb <= 3'b111;	end
		else if(x==43 && y==23) begin	rgb <= 3'b101;	end
		else if(x==44 && y==23) begin	rgb <= 3'b101;	end
		else if(x==5 && y==24) begin	rgb <= 3'b101;	end
		else if(x==6 && y==24) begin	rgb <= 3'b101;	end
		else if(x==7 && y==24) begin	rgb <= 3'b111;	end
		else if(x==8 && y==24) begin	rgb <= 3'b111;	end
		else if(x==9 && y==24) begin	rgb <= 3'b111;	end
		else if(x==10 && y==24) begin	rgb <= 3'b111;	end
		else if(x==11 && y==24) begin	rgb <= 3'b111;	end
		else if(x==12 && y==24) begin	rgb <= 3'b111;	end
		else if(x==13 && y==24) begin	rgb <= 3'b111;	end
		else if(x==14 && y==24) begin	rgb <= 3'b111;	end
		else if(x==15 && y==24) begin	rgb <= 3'b101;	end
		else if(x==16 && y==24) begin	rgb <= 3'b101;	end
		else if(x==17 && y==24) begin	rgb <= 3'b111;	end
		else if(x==18 && y==24) begin	rgb <= 3'b111;	end
		else if(x==19 && y==24) begin	rgb <= 3'b111;	end
		else if(x==20 && y==24) begin	rgb <= 3'b111;	end
		else if(x==21 && y==24) begin	rgb <= 3'b111;	end
		else if(x==22 && y==24) begin	rgb <= 3'b111;	end
		else if(x==23 && y==24) begin	rgb <= 3'b101;	end
		else if(x==24 && y==24) begin	rgb <= 3'b101;	end
		else if(x==25 && y==24) begin	rgb <= 3'b111;	end
		else if(x==26 && y==24) begin	rgb <= 3'b111;	end
		else if(x==27 && y==24) begin	rgb <= 3'b111;	end
		else if(x==28 && y==24) begin	rgb <= 3'b101;	end
		else if(x==29 && y==24) begin	rgb <= 3'b101;	end
		else if(x==30 && y==24) begin	rgb <= 3'b111;	end
		else if(x==31 && y==24) begin	rgb <= 3'b111;	end
		else if(x==32 && y==24) begin	rgb <= 3'b111;	end
		else if(x==33 && y==24) begin	rgb <= 3'b101;	end
		else if(x==34 && y==24) begin	rgb <= 3'b101;	end
		else if(x==35 && y==24) begin	rgb <= 3'b111;	end
		else if(x==36 && y==24) begin	rgb <= 3'b111;	end
		else if(x==37 && y==24) begin	rgb <= 3'b111;	end
		else if(x==38 && y==24) begin	rgb <= 3'b111;	end
		else if(x==39 && y==24) begin	rgb <= 3'b111;	end
		else if(x==40 && y==24) begin	rgb <= 3'b111;	end
		else if(x==41 && y==24) begin	rgb <= 3'b111;	end
		else if(x==42 && y==24) begin	rgb <= 3'b111;	end
		else if(x==43 && y==24) begin	rgb <= 3'b101;	end
		else if(x==44 && y==24) begin	rgb <= 3'b101;	end
		else if(x==2 && y==25) begin	rgb <= 3'b101;	end
		else if(x==3 && y==25) begin	rgb <= 3'b101;	end
		else if(x==4 && y==25) begin	rgb <= 3'b101;	end
		else if(x==5 && y==25) begin	rgb <= 3'b101;	end
		else if(x==6 && y==25) begin	rgb <= 3'b101;	end
		else if(x==7 && y==25) begin	rgb <= 3'b111;	end
		else if(x==8 && y==25) begin	rgb <= 3'b111;	end
		else if(x==9 && y==25) begin	rgb <= 3'b111;	end
		else if(x==10 && y==25) begin	rgb <= 3'b111;	end
		else if(x==11 && y==25) begin	rgb <= 3'b111;	end
		else if(x==12 && y==25) begin	rgb <= 3'b111;	end
		else if(x==13 && y==25) begin	rgb <= 3'b101;	end
		else if(x==14 && y==25) begin	rgb <= 3'b101;	end
		else if(x==15 && y==25) begin	rgb <= 3'b111;	end
		else if(x==16 && y==25) begin	rgb <= 3'b111;	end
		else if(x==17 && y==25) begin	rgb <= 3'b101;	end
		else if(x==20 && y==25) begin	rgb <= 3'b111;	end
		else if(x==21 && y==25) begin	rgb <= 3'b111;	end
		else if(x==22 && y==25) begin	rgb <= 3'b111;	end
		else if(x==23 && y==25) begin	rgb <= 3'b111;	end
		else if(x==24 && y==25) begin	rgb <= 3'b111;	end
		else if(x==25 && y==25) begin	rgb <= 3'b101;	end
		else if(x==26 && y==25) begin	rgb <= 3'b101;	end
		else if(x==27 && y==25) begin	rgb <= 3'b111;	end
		else if(x==28 && y==25) begin	rgb <= 3'b111;	end
		else if(x==29 && y==25) begin	rgb <= 3'b111;	end
		else if(x==32 && y==25) begin	rgb <= 3'b111;	end
		else if(x==33 && y==25) begin	rgb <= 3'b111;	end
		else if(x==34 && y==25) begin	rgb <= 3'b111;	end
		else if(x==35 && y==25) begin	rgb <= 3'b101;	end
		else if(x==36 && y==25) begin	rgb <= 3'b101;	end
		else if(x==37 && y==25) begin	rgb <= 3'b111;	end
		else if(x==38 && y==25) begin	rgb <= 3'b111;	end
		else if(x==39 && y==25) begin	rgb <= 3'b111;	end
		else if(x==40 && y==25) begin	rgb <= 3'b111;	end
		else if(x==41 && y==25) begin	rgb <= 3'b111;	end
		else if(x==42 && y==25) begin	rgb <= 3'b111;	end
		else if(x==43 && y==25) begin	rgb <= 3'b101;	end
		else if(x==44 && y==25) begin	rgb <= 3'b101;	end
		else if(x==45 && y==25) begin	rgb <= 3'b101;	end
		else if(x==46 && y==25) begin	rgb <= 3'b101;	end
		else if(x==2 && y==26) begin	rgb <= 3'b101;	end
		else if(x==3 && y==26) begin	rgb <= 3'b101;	end
		else if(x==4 && y==26) begin	rgb <= 3'b101;	end
		else if(x==5 && y==26) begin	rgb <= 3'b101;	end
		else if(x==6 && y==26) begin	rgb <= 3'b101;	end
		else if(x==7 && y==26) begin	rgb <= 3'b111;	end
		else if(x==8 && y==26) begin	rgb <= 3'b111;	end
		else if(x==9 && y==26) begin	rgb <= 3'b111;	end
		else if(x==10 && y==26) begin	rgb <= 3'b111;	end
		else if(x==11 && y==26) begin	rgb <= 3'b111;	end
		else if(x==12 && y==26) begin	rgb <= 3'b111;	end
		else if(x==13 && y==26) begin	rgb <= 3'b101;	end
		else if(x==14 && y==26) begin	rgb <= 3'b101;	end
		else if(x==15 && y==26) begin	rgb <= 3'b111;	end
		else if(x==16 && y==26) begin	rgb <= 3'b111;	end
		else if(x==17 && y==26) begin	rgb <= 3'b111;	end
		else if(x==20 && y==26) begin	rgb <= 3'b111;	end
		else if(x==21 && y==26) begin	rgb <= 3'b111;	end
		else if(x==22 && y==26) begin	rgb <= 3'b111;	end
		else if(x==23 && y==26) begin	rgb <= 3'b111;	end
		else if(x==24 && y==26) begin	rgb <= 3'b111;	end
		else if(x==25 && y==26) begin	rgb <= 3'b101;	end
		else if(x==26 && y==26) begin	rgb <= 3'b101;	end
		else if(x==27 && y==26) begin	rgb <= 3'b111;	end
		else if(x==28 && y==26) begin	rgb <= 3'b111;	end
		else if(x==29 && y==26) begin	rgb <= 3'b111;	end
		else if(x==32 && y==26) begin	rgb <= 3'b111;	end
		else if(x==33 && y==26) begin	rgb <= 3'b111;	end
		else if(x==34 && y==26) begin	rgb <= 3'b111;	end
		else if(x==35 && y==26) begin	rgb <= 3'b101;	end
		else if(x==36 && y==26) begin	rgb <= 3'b101;	end
		else if(x==37 && y==26) begin	rgb <= 3'b111;	end
		else if(x==38 && y==26) begin	rgb <= 3'b111;	end
		else if(x==39 && y==26) begin	rgb <= 3'b111;	end
		else if(x==40 && y==26) begin	rgb <= 3'b111;	end
		else if(x==41 && y==26) begin	rgb <= 3'b111;	end
		else if(x==42 && y==26) begin	rgb <= 3'b111;	end
		else if(x==43 && y==26) begin	rgb <= 3'b101;	end
		else if(x==44 && y==26) begin	rgb <= 3'b101;	end
		else if(x==45 && y==26) begin	rgb <= 3'b101;	end
		else if(x==46 && y==26) begin	rgb <= 3'b101;	end
		else if(x==1 && y==27) begin	rgb <= 3'b101;	end
		else if(x==2 && y==27) begin	rgb <= 3'b101;	end
		else if(x==3 && y==27) begin	rgb <= 3'b101;	end
		else if(x==4 && y==27) begin	rgb <= 3'b101;	end
		else if(x==7 && y==27) begin	rgb <= 3'b101;	end
		else if(x==8 && y==27) begin	rgb <= 3'b101;	end
		else if(x==9 && y==27) begin	rgb <= 3'b101;	end
		else if(x==10 && y==27) begin	rgb <= 3'b111;	end
		else if(x==11 && y==27) begin	rgb <= 3'b111;	end
		else if(x==12 && y==27) begin	rgb <= 3'b111;	end
		else if(x==13 && y==27) begin	rgb <= 3'b101;	end
		else if(x==14 && y==27) begin	rgb <= 3'b101;	end
		else if(x==15 && y==27) begin	rgb <= 3'b111;	end
		else if(x==16 && y==27) begin	rgb <= 3'b111;	end
		else if(x==17 && y==27) begin	rgb <= 3'b111;	end
		else if(x==18 && y==27) begin	rgb <= 3'b001;	end
		else if(x==19 && y==27) begin	rgb <= 3'b001;	end
		else if(x==20 && y==27) begin	rgb <= 3'b111;	end
		else if(x==21 && y==27) begin	rgb <= 3'b111;	end
		else if(x==22 && y==27) begin	rgb <= 3'b111;	end
		else if(x==23 && y==27) begin	rgb <= 3'b111;	end
		else if(x==24 && y==27) begin	rgb <= 3'b111;	end
		else if(x==25 && y==27) begin	rgb <= 3'b111;	end
		else if(x==26 && y==27) begin	rgb <= 3'b111;	end
		else if(x==27 && y==27) begin	rgb <= 3'b111;	end
		else if(x==28 && y==27) begin	rgb <= 3'b111;	end
		else if(x==29 && y==27) begin	rgb <= 3'b111;	end
		else if(x==30 && y==27) begin	rgb <= 3'b001;	end
		else if(x==31 && y==27) begin	rgb <= 3'b001;	end
		else if(x==32 && y==27) begin	rgb <= 3'b111;	end
		else if(x==33 && y==27) begin	rgb <= 3'b111;	end
		else if(x==34 && y==27) begin	rgb <= 3'b111;	end
		else if(x==35 && y==27) begin	rgb <= 3'b101;	end
		else if(x==36 && y==27) begin	rgb <= 3'b101;	end
		else if(x==37 && y==27) begin	rgb <= 3'b111;	end
		else if(x==38 && y==27) begin	rgb <= 3'b111;	end
		else if(x==39 && y==27) begin	rgb <= 3'b111;	end
		else if(x==40 && y==27) begin	rgb <= 3'b101;	end
		else if(x==41 && y==27) begin	rgb <= 3'b101;	end
		else if(x==45 && y==27) begin	rgb <= 3'b101;	end
		else if(x==46 && y==27) begin	rgb <= 3'b101;	end
		else if(x==47 && y==27) begin	rgb <= 3'b101;	end
		else if(x==48 && y==27) begin	rgb <= 3'b101;	end
		else if(x==49 && y==27) begin	rgb <= 3'b101;	end
		else if(x==1 && y==28) begin	rgb <= 3'b101;	end
		else if(x==2 && y==28) begin	rgb <= 3'b101;	end
		else if(x==3 && y==28) begin	rgb <= 3'b101;	end
		else if(x==4 && y==28) begin	rgb <= 3'b101;	end
		else if(x==7 && y==28) begin	rgb <= 3'b101;	end
		else if(x==8 && y==28) begin	rgb <= 3'b101;	end
		else if(x==9 && y==28) begin	rgb <= 3'b101;	end
		else if(x==10 && y==28) begin	rgb <= 3'b111;	end
		else if(x==11 && y==28) begin	rgb <= 3'b111;	end
		else if(x==12 && y==28) begin	rgb <= 3'b111;	end
		else if(x==13 && y==28) begin	rgb <= 3'b101;	end
		else if(x==14 && y==28) begin	rgb <= 3'b101;	end
		else if(x==15 && y==28) begin	rgb <= 3'b111;	end
		else if(x==16 && y==28) begin	rgb <= 3'b111;	end
		else if(x==17 && y==28) begin	rgb <= 3'b111;	end
		else if(x==18 && y==28) begin	rgb <= 3'b001;	end
		else if(x==19 && y==28) begin	rgb <= 3'b001;	end
		else if(x==20 && y==28) begin	rgb <= 3'b111;	end
		else if(x==21 && y==28) begin	rgb <= 3'b111;	end
		else if(x==22 && y==28) begin	rgb <= 3'b111;	end
		else if(x==23 && y==28) begin	rgb <= 3'b111;	end
		else if(x==24 && y==28) begin	rgb <= 3'b111;	end
		else if(x==25 && y==28) begin	rgb <= 3'b111;	end
		else if(x==26 && y==28) begin	rgb <= 3'b111;	end
		else if(x==27 && y==28) begin	rgb <= 3'b111;	end
		else if(x==28 && y==28) begin	rgb <= 3'b111;	end
		else if(x==29 && y==28) begin	rgb <= 3'b111;	end
		else if(x==30 && y==28) begin	rgb <= 3'b001;	end
		else if(x==31 && y==28) begin	rgb <= 3'b001;	end
		else if(x==32 && y==28) begin	rgb <= 3'b111;	end
		else if(x==33 && y==28) begin	rgb <= 3'b111;	end
		else if(x==34 && y==28) begin	rgb <= 3'b111;	end
		else if(x==35 && y==28) begin	rgb <= 3'b101;	end
		else if(x==36 && y==28) begin	rgb <= 3'b101;	end
		else if(x==37 && y==28) begin	rgb <= 3'b111;	end
		else if(x==38 && y==28) begin	rgb <= 3'b111;	end
		else if(x==39 && y==28) begin	rgb <= 3'b111;	end
		else if(x==40 && y==28) begin	rgb <= 3'b101;	end
		else if(x==41 && y==28) begin	rgb <= 3'b101;	end
		else if(x==45 && y==28) begin	rgb <= 3'b101;	end
		else if(x==46 && y==28) begin	rgb <= 3'b101;	end
		else if(x==47 && y==28) begin	rgb <= 3'b101;	end
		else if(x==48 && y==28) begin	rgb <= 3'b101;	end
		else if(x==49 && y==28) begin	rgb <= 3'b101;	end
		else if(x==1 && y==29) begin	rgb <= 3'b101;	end
		else if(x==2 && y==29) begin	rgb <= 3'b101;	end
		else if(x==3 && y==29) begin	rgb <= 3'b101;	end
		else if(x==4 && y==29) begin	rgb <= 3'b101;	end
		else if(x==7 && y==29) begin	rgb <= 3'b101;	end
		else if(x==8 && y==29) begin	rgb <= 3'b101;	end
		else if(x==9 && y==29) begin	rgb <= 3'b101;	end
		else if(x==10 && y==29) begin	rgb <= 3'b111;	end
		else if(x==11 && y==29) begin	rgb <= 3'b111;	end
		else if(x==12 && y==29) begin	rgb <= 3'b111;	end
		else if(x==13 && y==29) begin	rgb <= 3'b101;	end
		else if(x==14 && y==29) begin	rgb <= 3'b101;	end
		else if(x==15 && y==29) begin	rgb <= 3'b111;	end
		else if(x==16 && y==29) begin	rgb <= 3'b111;	end
		else if(x==17 && y==29) begin	rgb <= 3'b111;	end
		else if(x==18 && y==29) begin	rgb <= 3'b001;	end
		else if(x==19 && y==29) begin	rgb <= 3'b001;	end
		else if(x==20 && y==29) begin	rgb <= 3'b111;	end
		else if(x==21 && y==29) begin	rgb <= 3'b111;	end
		else if(x==22 && y==29) begin	rgb <= 3'b111;	end
		else if(x==23 && y==29) begin	rgb <= 3'b111;	end
		else if(x==24 && y==29) begin	rgb <= 3'b111;	end
		else if(x==25 && y==29) begin	rgb <= 3'b111;	end
		else if(x==26 && y==29) begin	rgb <= 3'b111;	end
		else if(x==27 && y==29) begin	rgb <= 3'b111;	end
		else if(x==28 && y==29) begin	rgb <= 3'b111;	end
		else if(x==29 && y==29) begin	rgb <= 3'b111;	end
		else if(x==30 && y==29) begin	rgb <= 3'b001;	end
		else if(x==31 && y==29) begin	rgb <= 3'b001;	end
		else if(x==32 && y==29) begin	rgb <= 3'b111;	end
		else if(x==33 && y==29) begin	rgb <= 3'b111;	end
		else if(x==34 && y==29) begin	rgb <= 3'b111;	end
		else if(x==35 && y==29) begin	rgb <= 3'b101;	end
		else if(x==36 && y==29) begin	rgb <= 3'b101;	end
		else if(x==37 && y==29) begin	rgb <= 3'b111;	end
		else if(x==38 && y==29) begin	rgb <= 3'b111;	end
		else if(x==39 && y==29) begin	rgb <= 3'b111;	end
		else if(x==40 && y==29) begin	rgb <= 3'b101;	end
		else if(x==41 && y==29) begin	rgb <= 3'b101;	end
		else if(x==45 && y==29) begin	rgb <= 3'b101;	end
		else if(x==46 && y==29) begin	rgb <= 3'b101;	end
		else if(x==47 && y==29) begin	rgb <= 3'b101;	end
		else if(x==48 && y==29) begin	rgb <= 3'b101;	end
		else if(x==49 && y==29) begin	rgb <= 3'b101;	end
		else if(x==7 && y==30) begin	rgb <= 3'b101;	end
		else if(x==8 && y==30) begin	rgb <= 3'b101;	end
		else if(x==9 && y==30) begin	rgb <= 3'b101;	end
		else if(x==10 && y==30) begin	rgb <= 3'b111;	end
		else if(x==11 && y==30) begin	rgb <= 3'b111;	end
		else if(x==12 && y==30) begin	rgb <= 3'b111;	end
		else if(x==13 && y==30) begin	rgb <= 3'b101;	end
		else if(x==14 && y==30) begin	rgb <= 3'b101;	end
		else if(x==15 && y==30) begin	rgb <= 3'b111;	end
		else if(x==16 && y==30) begin	rgb <= 3'b111;	end
		else if(x==17 && y==30) begin	rgb <= 3'b111;	end
		else if(x==18 && y==30) begin	rgb <= 3'b111;	end
		else if(x==19 && y==30) begin	rgb <= 3'b111;	end
		else if(x==20 && y==30) begin	rgb <= 3'b111;	end
		else if(x==21 && y==30) begin	rgb <= 3'b111;	end
		else if(x==22 && y==30) begin	rgb <= 3'b111;	end
		else if(x==23 && y==30) begin	rgb <= 3'b101;	end
		else if(x==24 && y==30) begin	rgb <= 3'b101;	end
		else if(x==25 && y==30) begin	rgb <= 3'b101;	end
		else if(x==26 && y==30) begin	rgb <= 3'b101;	end
		else if(x==27 && y==30) begin	rgb <= 3'b111;	end
		else if(x==28 && y==30) begin	rgb <= 3'b111;	end
		else if(x==29 && y==30) begin	rgb <= 3'b111;	end
		else if(x==30 && y==30) begin	rgb <= 3'b111;	end
		else if(x==31 && y==30) begin	rgb <= 3'b111;	end
		else if(x==32 && y==30) begin	rgb <= 3'b111;	end
		else if(x==33 && y==30) begin	rgb <= 3'b111;	end
		else if(x==34 && y==30) begin	rgb <= 3'b111;	end
		else if(x==35 && y==30) begin	rgb <= 3'b101;	end
		else if(x==36 && y==30) begin	rgb <= 3'b101;	end
		else if(x==37 && y==30) begin	rgb <= 3'b111;	end
		else if(x==38 && y==30) begin	rgb <= 3'b111;	end
		else if(x==39 && y==30) begin	rgb <= 3'b111;	end
		else if(x==40 && y==30) begin	rgb <= 3'b101;	end
		else if(x==41 && y==30) begin	rgb <= 3'b101;	end
		else if(x==7 && y==31) begin	rgb <= 3'b101;	end
		else if(x==8 && y==31) begin	rgb <= 3'b101;	end
		else if(x==9 && y==31) begin	rgb <= 3'b101;	end
		else if(x==10 && y==31) begin	rgb <= 3'b111;	end
		else if(x==11 && y==31) begin	rgb <= 3'b111;	end
		else if(x==12 && y==31) begin	rgb <= 3'b111;	end
		else if(x==13 && y==31) begin	rgb <= 3'b101;	end
		else if(x==14 && y==31) begin	rgb <= 3'b101;	end
		else if(x==15 && y==31) begin	rgb <= 3'b111;	end
		else if(x==16 && y==31) begin	rgb <= 3'b111;	end
		else if(x==17 && y==31) begin	rgb <= 3'b111;	end
		else if(x==18 && y==31) begin	rgb <= 3'b111;	end
		else if(x==19 && y==31) begin	rgb <= 3'b111;	end
		else if(x==20 && y==31) begin	rgb <= 3'b111;	end
		else if(x==21 && y==31) begin	rgb <= 3'b111;	end
		else if(x==22 && y==31) begin	rgb <= 3'b111;	end
		else if(x==23 && y==31) begin	rgb <= 3'b101;	end
		else if(x==24 && y==31) begin	rgb <= 3'b101;	end
		else if(x==25 && y==31) begin	rgb <= 3'b101;	end
		else if(x==26 && y==31) begin	rgb <= 3'b101;	end
		else if(x==27 && y==31) begin	rgb <= 3'b111;	end
		else if(x==28 && y==31) begin	rgb <= 3'b111;	end
		else if(x==29 && y==31) begin	rgb <= 3'b111;	end
		else if(x==30 && y==31) begin	rgb <= 3'b111;	end
		else if(x==31 && y==31) begin	rgb <= 3'b111;	end
		else if(x==32 && y==31) begin	rgb <= 3'b111;	end
		else if(x==33 && y==31) begin	rgb <= 3'b111;	end
		else if(x==34 && y==31) begin	rgb <= 3'b111;	end
		else if(x==35 && y==31) begin	rgb <= 3'b101;	end
		else if(x==36 && y==31) begin	rgb <= 3'b101;	end
		else if(x==37 && y==31) begin	rgb <= 3'b111;	end
		else if(x==38 && y==31) begin	rgb <= 3'b111;	end
		else if(x==39 && y==31) begin	rgb <= 3'b111;	end
		else if(x==40 && y==31) begin	rgb <= 3'b101;	end
		else if(x==41 && y==31) begin	rgb <= 3'b101;	end
		else if(x==42 && y==31) begin	rgb <= 3'b101;	end
		else if(x==10 && y==32) begin	rgb <= 3'b111;	end
		else if(x==11 && y==32) begin	rgb <= 3'b111;	end
		else if(x==12 && y==32) begin	rgb <= 3'b111;	end
		else if(x==13 && y==32) begin	rgb <= 3'b101;	end
		else if(x==14 && y==32) begin	rgb <= 3'b101;	end
		else if(x==15 && y==32) begin	rgb <= 3'b100;	end
		else if(x==16 && y==32) begin	rgb <= 3'b100;	end
		else if(x==17 && y==32) begin	rgb <= 3'b111;	end
		else if(x==18 && y==32) begin	rgb <= 3'b111;	end
		else if(x==19 && y==32) begin	rgb <= 3'b111;	end
		else if(x==20 && y==32) begin	rgb <= 3'b111;	end
		else if(x==21 && y==32) begin	rgb <= 3'b111;	end
		else if(x==22 && y==32) begin	rgb <= 3'b111;	end
		else if(x==23 && y==32) begin	rgb <= 3'b111;	end
		else if(x==24 && y==32) begin	rgb <= 3'b111;	end
		else if(x==25 && y==32) begin	rgb <= 3'b111;	end
		else if(x==26 && y==32) begin	rgb <= 3'b111;	end
		else if(x==27 && y==32) begin	rgb <= 3'b111;	end
		else if(x==28 && y==32) begin	rgb <= 3'b111;	end
		else if(x==29 && y==32) begin	rgb <= 3'b111;	end
		else if(x==30 && y==32) begin	rgb <= 3'b111;	end
		else if(x==31 && y==32) begin	rgb <= 3'b111;	end
		else if(x==32 && y==32) begin	rgb <= 3'b111;	end
		else if(x==33 && y==32) begin	rgb <= 3'b100;	end
		else if(x==34 && y==32) begin	rgb <= 3'b100;	end
		else if(x==35 && y==32) begin	rgb <= 3'b101;	end
		else if(x==36 && y==32) begin	rgb <= 3'b101;	end
		else if(x==37 && y==32) begin	rgb <= 3'b111;	end
		else if(x==38 && y==32) begin	rgb <= 3'b111;	end
		else if(x==39 && y==32) begin	rgb <= 3'b111;	end
		else if(x==10 && y==33) begin	rgb <= 3'b111;	end
		else if(x==11 && y==33) begin	rgb <= 3'b111;	end
		else if(x==12 && y==33) begin	rgb <= 3'b111;	end
		else if(x==13 && y==33) begin	rgb <= 3'b101;	end
		else if(x==14 && y==33) begin	rgb <= 3'b101;	end
		else if(x==15 && y==33) begin	rgb <= 3'b100;	end
		else if(x==16 && y==33) begin	rgb <= 3'b100;	end
		else if(x==17 && y==33) begin	rgb <= 3'b111;	end
		else if(x==18 && y==33) begin	rgb <= 3'b111;	end
		else if(x==19 && y==33) begin	rgb <= 3'b111;	end
		else if(x==20 && y==33) begin	rgb <= 3'b111;	end
		else if(x==21 && y==33) begin	rgb <= 3'b111;	end
		else if(x==22 && y==33) begin	rgb <= 3'b111;	end
		else if(x==23 && y==33) begin	rgb <= 3'b111;	end
		else if(x==24 && y==33) begin	rgb <= 3'b111;	end
		else if(x==25 && y==33) begin	rgb <= 3'b111;	end
		else if(x==26 && y==33) begin	rgb <= 3'b111;	end
		else if(x==27 && y==33) begin	rgb <= 3'b111;	end
		else if(x==28 && y==33) begin	rgb <= 3'b111;	end
		else if(x==29 && y==33) begin	rgb <= 3'b111;	end
		else if(x==30 && y==33) begin	rgb <= 3'b111;	end
		else if(x==31 && y==33) begin	rgb <= 3'b111;	end
		else if(x==32 && y==33) begin	rgb <= 3'b111;	end
		else if(x==33 && y==33) begin	rgb <= 3'b100;	end
		else if(x==34 && y==33) begin	rgb <= 3'b100;	end
		else if(x==35 && y==33) begin	rgb <= 3'b101;	end
		else if(x==36 && y==33) begin	rgb <= 3'b101;	end
		else if(x==37 && y==33) begin	rgb <= 3'b111;	end
		else if(x==38 && y==33) begin	rgb <= 3'b111;	end
		else if(x==39 && y==33) begin	rgb <= 3'b111;	end
		else if(x==7 && y==34) begin	rgb <= 3'b101;	end
		else if(x==8 && y==34) begin	rgb <= 3'b101;	end
		else if(x==9 && y==34) begin	rgb <= 3'b101;	end
		else if(x==10 && y==34) begin	rgb <= 3'b111;	end
		else if(x==11 && y==34) begin	rgb <= 3'b111;	end
		else if(x==12 && y==34) begin	rgb <= 3'b111;	end
		else if(x==13 && y==34) begin	rgb <= 3'b111;	end
		else if(x==14 && y==34) begin	rgb <= 3'b111;	end
		else if(x==15 && y==34) begin	rgb <= 3'b100;	end
		else if(x==16 && y==34) begin	rgb <= 3'b100;	end
		else if(x==17 && y==34) begin	rgb <= 3'b100;	end
		else if(x==18 && y==34) begin	rgb <= 3'b100;	end
		else if(x==19 && y==34) begin	rgb <= 3'b100;	end
		else if(x==20 && y==34) begin	rgb <= 3'b100;	end
		else if(x==21 && y==34) begin	rgb <= 3'b100;	end
		else if(x==27 && y==34) begin	rgb <= 3'b100;	end
		else if(x==28 && y==34) begin	rgb <= 3'b100;	end
		else if(x==29 && y==34) begin	rgb <= 3'b100;	end
		else if(x==30 && y==34) begin	rgb <= 3'b100;	end
		else if(x==31 && y==34) begin	rgb <= 3'b100;	end
		else if(x==32 && y==34) begin	rgb <= 3'b100;	end
		else if(x==33 && y==34) begin	rgb <= 3'b100;	end
		else if(x==34 && y==34) begin	rgb <= 3'b100;	end
		else if(x==35 && y==34) begin	rgb <= 3'b111;	end
		else if(x==36 && y==34) begin	rgb <= 3'b111;	end
		else if(x==37 && y==34) begin	rgb <= 3'b111;	end
		else if(x==38 && y==34) begin	rgb <= 3'b111;	end
		else if(x==39 && y==34) begin	rgb <= 3'b111;	end
		else if(x==40 && y==34) begin	rgb <= 3'b101;	end
		else if(x==41 && y==34) begin	rgb <= 3'b101;	end
		else if(x==7 && y==35) begin	rgb <= 3'b101;	end
		else if(x==8 && y==35) begin	rgb <= 3'b101;	end
		else if(x==9 && y==35) begin	rgb <= 3'b101;	end
		else if(x==10 && y==35) begin	rgb <= 3'b111;	end
		else if(x==11 && y==35) begin	rgb <= 3'b111;	end
		else if(x==12 && y==35) begin	rgb <= 3'b111;	end
		else if(x==13 && y==35) begin	rgb <= 3'b111;	end
		else if(x==14 && y==35) begin	rgb <= 3'b111;	end
		else if(x==15 && y==35) begin	rgb <= 3'b100;	end
		else if(x==16 && y==35) begin	rgb <= 3'b100;	end
		else if(x==17 && y==35) begin	rgb <= 3'b100;	end
		else if(x==18 && y==35) begin	rgb <= 3'b100;	end
		else if(x==19 && y==35) begin	rgb <= 3'b100;	end
		else if(x==20 && y==35) begin	rgb <= 3'b100;	end
		else if(x==21 && y==35) begin	rgb <= 3'b100;	end
		else if(x==27 && y==35) begin	rgb <= 3'b100;	end
		else if(x==28 && y==35) begin	rgb <= 3'b100;	end
		else if(x==29 && y==35) begin	rgb <= 3'b100;	end
		else if(x==30 && y==35) begin	rgb <= 3'b100;	end
		else if(x==31 && y==35) begin	rgb <= 3'b100;	end
		else if(x==32 && y==35) begin	rgb <= 3'b100;	end
		else if(x==33 && y==35) begin	rgb <= 3'b100;	end
		else if(x==34 && y==35) begin	rgb <= 3'b100;	end
		else if(x==35 && y==35) begin	rgb <= 3'b111;	end
		else if(x==36 && y==35) begin	rgb <= 3'b111;	end
		else if(x==37 && y==35) begin	rgb <= 3'b111;	end
		else if(x==38 && y==35) begin	rgb <= 3'b111;	end
		else if(x==39 && y==35) begin	rgb <= 3'b111;	end
		else if(x==40 && y==35) begin	rgb <= 3'b101;	end
		else if(x==41 && y==35) begin	rgb <= 3'b101;	end
		else if(x==7 && y==36) begin	rgb <= 3'b101;	end
		else if(x==8 && y==36) begin	rgb <= 3'b101;	end
		else if(x==9 && y==36) begin	rgb <= 3'b101;	end
		else if(x==10 && y==36) begin	rgb <= 3'b111;	end
		else if(x==11 && y==36) begin	rgb <= 3'b111;	end
		else if(x==12 && y==36) begin	rgb <= 3'b111;	end
		else if(x==13 && y==36) begin	rgb <= 3'b111;	end
		else if(x==14 && y==36) begin	rgb <= 3'b111;	end
		else if(x==15 && y==36) begin	rgb <= 3'b100;	end
		else if(x==16 && y==36) begin	rgb <= 3'b100;	end
		else if(x==17 && y==36) begin	rgb <= 3'b100;	end
		else if(x==18 && y==36) begin	rgb <= 3'b100;	end
		else if(x==19 && y==36) begin	rgb <= 3'b100;	end
		else if(x==22 && y==36) begin	rgb <= 3'b111;	end
		else if(x==23 && y==36) begin	rgb <= 3'b111;	end
		else if(x==24 && y==36) begin	rgb <= 3'b111;	end
		else if(x==25 && y==36) begin	rgb <= 3'b111;	end
		else if(x==26 && y==36) begin	rgb <= 3'b111;	end
		else if(x==30 && y==36) begin	rgb <= 3'b100;	end
		else if(x==31 && y==36) begin	rgb <= 3'b100;	end
		else if(x==32 && y==36) begin	rgb <= 3'b100;	end
		else if(x==33 && y==36) begin	rgb <= 3'b100;	end
		else if(x==34 && y==36) begin	rgb <= 3'b100;	end
		else if(x==35 && y==36) begin	rgb <= 3'b111;	end
		else if(x==36 && y==36) begin	rgb <= 3'b111;	end
		else if(x==37 && y==36) begin	rgb <= 3'b111;	end
		else if(x==38 && y==36) begin	rgb <= 3'b111;	end
		else if(x==39 && y==36) begin	rgb <= 3'b111;	end
		else if(x==40 && y==36) begin	rgb <= 3'b101;	end
		else if(x==41 && y==36) begin	rgb <= 3'b101;	end
		else if(x==7 && y==37) begin	rgb <= 3'b101;	end
		else if(x==8 && y==37) begin	rgb <= 3'b101;	end
		else if(x==9 && y==37) begin	rgb <= 3'b101;	end
		else if(x==10 && y==37) begin	rgb <= 3'b111;	end
		else if(x==11 && y==37) begin	rgb <= 3'b111;	end
		else if(x==12 && y==37) begin	rgb <= 3'b111;	end
		else if(x==13 && y==37) begin	rgb <= 3'b111;	end
		else if(x==14 && y==37) begin	rgb <= 3'b111;	end
		else if(x==15 && y==37) begin	rgb <= 3'b100;	end
		else if(x==16 && y==37) begin	rgb <= 3'b100;	end
		else if(x==17 && y==37) begin	rgb <= 3'b100;	end
		else if(x==18 && y==37) begin	rgb <= 3'b100;	end
		else if(x==19 && y==37) begin	rgb <= 3'b100;	end
		else if(x==22 && y==37) begin	rgb <= 3'b111;	end
		else if(x==23 && y==37) begin	rgb <= 3'b111;	end
		else if(x==24 && y==37) begin	rgb <= 3'b111;	end
		else if(x==25 && y==37) begin	rgb <= 3'b111;	end
		else if(x==26 && y==37) begin	rgb <= 3'b111;	end
		else if(x==30 && y==37) begin	rgb <= 3'b100;	end
		else if(x==31 && y==37) begin	rgb <= 3'b100;	end
		else if(x==32 && y==37) begin	rgb <= 3'b100;	end
		else if(x==33 && y==37) begin	rgb <= 3'b100;	end
		else if(x==34 && y==37) begin	rgb <= 3'b100;	end
		else if(x==35 && y==37) begin	rgb <= 3'b111;	end
		else if(x==36 && y==37) begin	rgb <= 3'b111;	end
		else if(x==37 && y==37) begin	rgb <= 3'b111;	end
		else if(x==38 && y==37) begin	rgb <= 3'b111;	end
		else if(x==39 && y==37) begin	rgb <= 3'b111;	end
		else if(x==40 && y==37) begin	rgb <= 3'b101;	end
		else if(x==41 && y==37) begin	rgb <= 3'b101;	end
		else if(x==7 && y==38) begin	rgb <= 3'b101;	end
		else if(x==8 && y==38) begin	rgb <= 3'b101;	end
		else if(x==9 && y==38) begin	rgb <= 3'b101;	end
		else if(x==10 && y==38) begin	rgb <= 3'b111;	end
		else if(x==11 && y==38) begin	rgb <= 3'b111;	end
		else if(x==12 && y==38) begin	rgb <= 3'b111;	end
		else if(x==13 && y==38) begin	rgb <= 3'b111;	end
		else if(x==14 && y==38) begin	rgb <= 3'b111;	end
		else if(x==15 && y==38) begin	rgb <= 3'b100;	end
		else if(x==16 && y==38) begin	rgb <= 3'b100;	end
		else if(x==17 && y==38) begin	rgb <= 3'b100;	end
		else if(x==18 && y==38) begin	rgb <= 3'b100;	end
		else if(x==19 && y==38) begin	rgb <= 3'b100;	end
		else if(x==22 && y==38) begin	rgb <= 3'b100;	end
		else if(x==23 && y==38) begin	rgb <= 3'b111;	end
		else if(x==24 && y==38) begin	rgb <= 3'b111;	end
		else if(x==25 && y==38) begin	rgb <= 3'b111;	end
		else if(x==26 && y==38) begin	rgb <= 3'b111;	end
		else if(x==30 && y==38) begin	rgb <= 3'b100;	end
		else if(x==31 && y==38) begin	rgb <= 3'b100;	end
		else if(x==32 && y==38) begin	rgb <= 3'b100;	end
		else if(x==33 && y==38) begin	rgb <= 3'b100;	end
		else if(x==34 && y==38) begin	rgb <= 3'b100;	end
		else if(x==35 && y==38) begin	rgb <= 3'b111;	end
		else if(x==36 && y==38) begin	rgb <= 3'b111;	end
		else if(x==37 && y==38) begin	rgb <= 3'b111;	end
		else if(x==38 && y==38) begin	rgb <= 3'b111;	end
		else if(x==39 && y==38) begin	rgb <= 3'b111;	end
		else if(x==40 && y==38) begin	rgb <= 3'b101;	end
		else if(x==41 && y==38) begin	rgb <= 3'b101;	end
		else if(x==10 && y==39) begin	rgb <= 3'b111;	end
		else if(x==11 && y==39) begin	rgb <= 3'b111;	end
		else if(x==12 && y==39) begin	rgb <= 3'b111;	end
		else if(x==13 && y==39) begin	rgb <= 3'b101;	end
		else if(x==14 && y==39) begin	rgb <= 3'b101;	end
		else if(x==15 && y==39) begin	rgb <= 3'b100;	end
		else if(x==16 && y==39) begin	rgb <= 3'b100;	end
		else if(x==33 && y==39) begin	rgb <= 3'b100;	end
		else if(x==34 && y==39) begin	rgb <= 3'b100;	end
		else if(x==35 && y==39) begin	rgb <= 3'b101;	end
		else if(x==36 && y==39) begin	rgb <= 3'b101;	end
		else if(x==37 && y==39) begin	rgb <= 3'b111;	end
		else if(x==38 && y==39) begin	rgb <= 3'b111;	end
		else if(x==39 && y==39) begin	rgb <= 3'b111;	end
		else if(x==10 && y==40) begin	rgb <= 3'b111;	end
		else if(x==11 && y==40) begin	rgb <= 3'b111;	end
		else if(x==12 && y==40) begin	rgb <= 3'b111;	end
		else if(x==13 && y==40) begin	rgb <= 3'b101;	end
		else if(x==14 && y==40) begin	rgb <= 3'b101;	end
		else if(x==15 && y==40) begin	rgb <= 3'b100;	end
		else if(x==16 && y==40) begin	rgb <= 3'b100;	end
		else if(x==33 && y==40) begin	rgb <= 3'b100;	end
		else if(x==34 && y==40) begin	rgb <= 3'b100;	end
		else if(x==35 && y==40) begin	rgb <= 3'b101;	end
		else if(x==36 && y==40) begin	rgb <= 3'b101;	end
		else if(x==37 && y==40) begin	rgb <= 3'b111;	end
		else if(x==38 && y==40) begin	rgb <= 3'b111;	end
		else if(x==39 && y==40) begin	rgb <= 3'b111;	end
		else if(x==10 && y==41) begin	rgb <= 3'b111;	end
		else if(x==11 && y==41) begin	rgb <= 3'b111;	end
		else if(x==12 && y==41) begin	rgb <= 3'b111;	end
		else if(x==13 && y==41) begin	rgb <= 3'b101;	end
		else if(x==14 && y==41) begin	rgb <= 3'b101;	end
		else if(x==15 && y==41) begin	rgb <= 3'b111;	end
		else if(x==16 && y==41) begin	rgb <= 3'b111;	end
		else if(x==17 && y==41) begin	rgb <= 3'b111;	end
		else if(x==18 && y==41) begin	rgb <= 3'b100;	end
		else if(x==19 && y==41) begin	rgb <= 3'b100;	end
		else if(x==22 && y==41) begin	rgb <= 3'b101;	end
		else if(x==23 && y==41) begin	rgb <= 3'b101;	end
		else if(x==24 && y==41) begin	rgb <= 3'b101;	end
		else if(x==25 && y==41) begin	rgb <= 3'b101;	end
		else if(x==26 && y==41) begin	rgb <= 3'b101;	end
		else if(x==27 && y==41) begin	rgb <= 3'b101;	end
		else if(x==30 && y==41) begin	rgb <= 3'b100;	end
		else if(x==31 && y==41) begin	rgb <= 3'b100;	end
		else if(x==32 && y==41) begin	rgb <= 3'b111;	end
		else if(x==33 && y==41) begin	rgb <= 3'b111;	end
		else if(x==34 && y==41) begin	rgb <= 3'b111;	end
		else if(x==35 && y==41) begin	rgb <= 3'b101;	end
		else if(x==36 && y==41) begin	rgb <= 3'b101;	end
		else if(x==37 && y==41) begin	rgb <= 3'b111;	end
		else if(x==38 && y==41) begin	rgb <= 3'b111;	end
		else if(x==39 && y==41) begin	rgb <= 3'b111;	end
		else if(x==10 && y==42) begin	rgb <= 3'b111;	end
		else if(x==11 && y==42) begin	rgb <= 3'b111;	end
		else if(x==12 && y==42) begin	rgb <= 3'b111;	end
		else if(x==13 && y==42) begin	rgb <= 3'b101;	end
		else if(x==14 && y==42) begin	rgb <= 3'b101;	end
		else if(x==15 && y==42) begin	rgb <= 3'b111;	end
		else if(x==16 && y==42) begin	rgb <= 3'b111;	end
		else if(x==17 && y==42) begin	rgb <= 3'b111;	end
		else if(x==18 && y==42) begin	rgb <= 3'b100;	end
		else if(x==19 && y==42) begin	rgb <= 3'b100;	end
		else if(x==22 && y==42) begin	rgb <= 3'b101;	end
		else if(x==23 && y==42) begin	rgb <= 3'b101;	end
		else if(x==24 && y==42) begin	rgb <= 3'b101;	end
		else if(x==25 && y==42) begin	rgb <= 3'b101;	end
		else if(x==26 && y==42) begin	rgb <= 3'b101;	end
		else if(x==27 && y==42) begin	rgb <= 3'b101;	end
		else if(x==30 && y==42) begin	rgb <= 3'b100;	end
		else if(x==31 && y==42) begin	rgb <= 3'b100;	end
		else if(x==32 && y==42) begin	rgb <= 3'b111;	end
		else if(x==33 && y==42) begin	rgb <= 3'b111;	end
		else if(x==34 && y==42) begin	rgb <= 3'b111;	end
		else if(x==35 && y==42) begin	rgb <= 3'b101;	end
		else if(x==36 && y==42) begin	rgb <= 3'b101;	end
		else if(x==37 && y==42) begin	rgb <= 3'b111;	end
		else if(x==38 && y==42) begin	rgb <= 3'b111;	end
		else if(x==39 && y==42) begin	rgb <= 3'b111;	end
		else if(x==10 && y==43) begin	rgb <= 3'b111;	end
		else if(x==11 && y==43) begin	rgb <= 3'b111;	end
		else if(x==12 && y==43) begin	rgb <= 3'b111;	end
		else if(x==13 && y==43) begin	rgb <= 3'b101;	end
		else if(x==14 && y==43) begin	rgb <= 3'b101;	end
		else if(x==15 && y==43) begin	rgb <= 3'b100;	end
		else if(x==16 && y==43) begin	rgb <= 3'b100;	end
		else if(x==17 && y==43) begin	rgb <= 3'b101;	end
		else if(x==18 && y==43) begin	rgb <= 3'b101;	end
		else if(x==19 && y==43) begin	rgb <= 3'b101;	end
		else if(x==20 && y==43) begin	rgb <= 3'b101;	end
		else if(x==21 && y==43) begin	rgb <= 3'b101;	end
		else if(x==22 && y==43) begin	rgb <= 3'b101;	end
		else if(x==23 && y==43) begin	rgb <= 3'b101;	end
		else if(x==24 && y==43) begin	rgb <= 3'b101;	end
		else if(x==25 && y==43) begin	rgb <= 3'b101;	end
		else if(x==26 && y==43) begin	rgb <= 3'b101;	end
		else if(x==27 && y==43) begin	rgb <= 3'b101;	end
		else if(x==28 && y==43) begin	rgb <= 3'b101;	end
		else if(x==29 && y==43) begin	rgb <= 3'b101;	end
		else if(x==30 && y==43) begin	rgb <= 3'b101;	end
		else if(x==31 && y==43) begin	rgb <= 3'b101;	end
		else if(x==32 && y==43) begin	rgb <= 3'b101;	end
		else if(x==33 && y==43) begin	rgb <= 3'b100;	end
		else if(x==34 && y==43) begin	rgb <= 3'b100;	end
		else if(x==35 && y==43) begin	rgb <= 3'b101;	end
		else if(x==36 && y==43) begin	rgb <= 3'b101;	end
		else if(x==37 && y==43) begin	rgb <= 3'b111;	end
		else if(x==38 && y==43) begin	rgb <= 3'b111;	end
		else if(x==39 && y==43) begin	rgb <= 3'b111;	end
		else if(x==10 && y==44) begin	rgb <= 3'b111;	end
		else if(x==11 && y==44) begin	rgb <= 3'b111;	end
		else if(x==12 && y==44) begin	rgb <= 3'b111;	end
		else if(x==13 && y==44) begin	rgb <= 3'b101;	end
		else if(x==14 && y==44) begin	rgb <= 3'b101;	end
		else if(x==15 && y==44) begin	rgb <= 3'b100;	end
		else if(x==16 && y==44) begin	rgb <= 3'b100;	end
		else if(x==17 && y==44) begin	rgb <= 3'b101;	end
		else if(x==18 && y==44) begin	rgb <= 3'b101;	end
		else if(x==19 && y==44) begin	rgb <= 3'b101;	end
		else if(x==20 && y==44) begin	rgb <= 3'b101;	end
		else if(x==21 && y==44) begin	rgb <= 3'b101;	end
		else if(x==22 && y==44) begin	rgb <= 3'b101;	end
		else if(x==23 && y==44) begin	rgb <= 3'b101;	end
		else if(x==24 && y==44) begin	rgb <= 3'b101;	end
		else if(x==25 && y==44) begin	rgb <= 3'b101;	end
		else if(x==26 && y==44) begin	rgb <= 3'b101;	end
		else if(x==27 && y==44) begin	rgb <= 3'b101;	end
		else if(x==28 && y==44) begin	rgb <= 3'b101;	end
		else if(x==29 && y==44) begin	rgb <= 3'b101;	end
		else if(x==30 && y==44) begin	rgb <= 3'b101;	end
		else if(x==31 && y==44) begin	rgb <= 3'b101;	end
		else if(x==32 && y==44) begin	rgb <= 3'b101;	end
		else if(x==33 && y==44) begin	rgb <= 3'b100;	end
		else if(x==34 && y==44) begin	rgb <= 3'b100;	end
		else if(x==35 && y==44) begin	rgb <= 3'b101;	end
		else if(x==36 && y==44) begin	rgb <= 3'b101;	end
		else if(x==37 && y==44) begin	rgb <= 3'b111;	end
		else if(x==38 && y==44) begin	rgb <= 3'b111;	end
		else if(x==39 && y==44) begin	rgb <= 3'b111;	end
		else if(x==10 && y==45) begin	rgb <= 3'b101;	end
		else if(x==11 && y==45) begin	rgb <= 3'b101;	end
		else if(x==15 && y==45) begin	rgb <= 3'b100;	end
		else if(x==16 && y==45) begin	rgb <= 3'b100;	end
		else if(x==17 && y==45) begin	rgb <= 3'b100;	end
		else if(x==18 && y==45) begin	rgb <= 3'b100;	end
		else if(x==19 && y==45) begin	rgb <= 3'b100;	end
		else if(x==20 && y==45) begin	rgb <= 3'b111;	end
		else if(x==21 && y==45) begin	rgb <= 3'b111;	end
		else if(x==22 && y==45) begin	rgb <= 3'b111;	end
		else if(x==23 && y==45) begin	rgb <= 3'b100;	end
		else if(x==24 && y==45) begin	rgb <= 3'b100;	end
		else if(x==25 && y==45) begin	rgb <= 3'b100;	end
		else if(x==26 && y==45) begin	rgb <= 3'b100;	end
		else if(x==27 && y==45) begin	rgb <= 3'b111;	end
		else if(x==28 && y==45) begin	rgb <= 3'b111;	end
		else if(x==29 && y==45) begin	rgb <= 3'b111;	end
		else if(x==30 && y==45) begin	rgb <= 3'b100;	end
		else if(x==31 && y==45) begin	rgb <= 3'b100;	end
		else if(x==32 && y==45) begin	rgb <= 3'b100;	end
		else if(x==33 && y==45) begin	rgb <= 3'b100;	end
		else if(x==34 && y==45) begin	rgb <= 3'b100;	end
		else if(x==37 && y==45) begin	rgb <= 3'b101;	end
		else if(x==38 && y==45) begin	rgb <= 3'b101;	end
		else if(x==39 && y==45) begin	rgb <= 3'b101;	end
		else if(x==10 && y==46) begin	rgb <= 3'b101;	end
		else if(x==11 && y==46) begin	rgb <= 3'b101;	end
		else if(x==15 && y==46) begin	rgb <= 3'b100;	end
		else if(x==16 && y==46) begin	rgb <= 3'b100;	end
		else if(x==17 && y==46) begin	rgb <= 3'b100;	end
		else if(x==18 && y==46) begin	rgb <= 3'b100;	end
		else if(x==19 && y==46) begin	rgb <= 3'b100;	end
		else if(x==20 && y==46) begin	rgb <= 3'b111;	end
		else if(x==21 && y==46) begin	rgb <= 3'b111;	end
		else if(x==22 && y==46) begin	rgb <= 3'b111;	end
		else if(x==23 && y==46) begin	rgb <= 3'b100;	end
		else if(x==24 && y==46) begin	rgb <= 3'b100;	end
		else if(x==25 && y==46) begin	rgb <= 3'b100;	end
		else if(x==26 && y==46) begin	rgb <= 3'b100;	end
		else if(x==27 && y==46) begin	rgb <= 3'b111;	end
		else if(x==28 && y==46) begin	rgb <= 3'b111;	end
		else if(x==29 && y==46) begin	rgb <= 3'b111;	end
		else if(x==30 && y==46) begin	rgb <= 3'b100;	end
		else if(x==31 && y==46) begin	rgb <= 3'b100;	end
		else if(x==32 && y==46) begin	rgb <= 3'b100;	end
		else if(x==33 && y==46) begin	rgb <= 3'b100;	end
		else if(x==34 && y==46) begin	rgb <= 3'b100;	end
		else if(x==37 && y==46) begin	rgb <= 3'b101;	end
		else if(x==38 && y==46) begin	rgb <= 3'b101;	end
		else if(x==39 && y==46) begin	rgb <= 3'b101;	end
		else if(x==10 && y==47) begin	rgb <= 3'b101;	end
		else if(x==11 && y==47) begin	rgb <= 3'b101;	end
		else if(x==15 && y==47) begin	rgb <= 3'b100;	end
		else if(x==16 && y==47) begin	rgb <= 3'b100;	end
		else if(x==17 && y==47) begin	rgb <= 3'b100;	end
		else if(x==18 && y==47) begin	rgb <= 3'b100;	end
		else if(x==19 && y==47) begin	rgb <= 3'b100;	end
		else if(x==20 && y==47) begin	rgb <= 3'b111;	end
		else if(x==21 && y==47) begin	rgb <= 3'b111;	end
		else if(x==22 && y==47) begin	rgb <= 3'b111;	end
		else if(x==23 && y==47) begin	rgb <= 3'b100;	end
		else if(x==24 && y==47) begin	rgb <= 3'b100;	end
		else if(x==25 && y==47) begin	rgb <= 3'b100;	end
		else if(x==26 && y==47) begin	rgb <= 3'b100;	end
		else if(x==27 && y==47) begin	rgb <= 3'b111;	end
		else if(x==28 && y==47) begin	rgb <= 3'b111;	end
		else if(x==29 && y==47) begin	rgb <= 3'b111;	end
		else if(x==30 && y==47) begin	rgb <= 3'b100;	end
		else if(x==31 && y==47) begin	rgb <= 3'b100;	end
		else if(x==32 && y==47) begin	rgb <= 3'b100;	end
		else if(x==33 && y==47) begin	rgb <= 3'b100;	end
		else if(x==34 && y==47) begin	rgb <= 3'b100;	end
		else if(x==37 && y==47) begin	rgb <= 3'b101;	end
		else if(x==38 && y==47) begin	rgb <= 3'b101;	end
		else if(x==39 && y==47) begin	rgb <= 3'b101;	end
		else if(x==20 && y==48) begin	rgb <= 3'b111;	end
		else if(x==21 && y==48) begin	rgb <= 3'b111;	end
		else if(x==27 && y==48) begin	rgb <= 3'b111;	end
		else if(x==28 && y==48) begin	rgb <= 3'b111;	end
		else if(x==29 && y==48) begin	rgb <= 3'b111;	end
		else if(x==20 && y==49) begin	rgb <= 3'b111;	end
		else if(x==21 && y==49) begin	rgb <= 3'b111;	end
		else if(x==22 && y==49) begin	rgb <= 3'b111;	end
		else if(x==27 && y==49) begin	rgb <= 3'b111;	end
		else if(x==28 && y==49) begin	rgb <= 3'b111;	end
		else if(x==29 && y==49) begin	rgb <= 3'b111;	end
		else begin rgb <= 3'b000; end// Width: 50, Height: 50 From: C:/Users/ITPCC/Desktop/vocaloid-50.png
	end
endmodule